module mult_512_part (
    input wire clk,
    input wire CE,
    input wire rst,

    input wire [255 : 0] mult_part_in0,
    input wire [255 : 0] mult_part_in1,

    output reg [511 : 0] mult_part_out00,
    output reg [511 : 0] mult_part_out01,
    output reg [511 : 0] mult_part_out02,
    output reg [511 : 0] mult_part_out03,
    output reg [511 : 0] mult_part_out04,
    output reg [511 : 0] mult_part_out05,
    output reg [511 : 0] mult_part_out06,
    output reg [511 : 0] mult_part_out07,
    output reg [511 : 0] mult_part_out08,
    output reg [511 : 0] mult_part_out09,
    output reg [511 : 0] mult_part_out10,
    output reg [511 : 0] mult_part_out11,
    output reg [511 : 0] mult_part_out12,
    output reg [511 : 0] mult_part_out13,
    output reg [511 : 0] mult_part_out14,
    output reg [511 : 0] mult_part_out15,
    output reg [511 : 0] mult_part_out16,
    output reg [511 : 0] mult_part_out17,
    output reg [511 : 0] mult_part_out18,
    output reg [511 : 0] mult_part_out19,
    output reg [511 : 0] mult_part_out20,
    output reg [511 : 0] mult_part_out21,
    output reg [511 : 0] mult_part_out22,
    output reg [511 : 0] mult_part_out23,
    output reg [511 : 0] mult_part_out24,
    output reg [511 : 0] mult_part_out25
    );


wire [42 : 0] P_0_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_0 (
  .P(P_0_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_1 (
  .P(P_0_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_2 (
  .P(P_0_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_3 (
  .P(P_0_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_4 (
  .P(P_0_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_5 (
  .P(P_0_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_6 (
  .P(P_0_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_7 (
  .P(P_0_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_8 (
  .P(P_0_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_0_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_9 (
  .P(P_0_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_0_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_0_10 (
  .P(P_0_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[16:0]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_0 (
  .P(P_1_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_1 (
  .P(P_1_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_2 (
  .P(P_1_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_3 (
  .P(P_1_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_4 (
  .P(P_1_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_5 (
  .P(P_1_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_6 (
  .P(P_1_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_7 (
  .P(P_1_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_8 (
  .P(P_1_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_1_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_9 (
  .P(P_1_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_1_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_1_10 (
  .P(P_1_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[33:17]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_0 (
  .P(P_2_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_1 (
  .P(P_2_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_2 (
  .P(P_2_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_3 (
  .P(P_2_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_4 (
  .P(P_2_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_5 (
  .P(P_2_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_6 (
  .P(P_2_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_7 (
  .P(P_2_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_8 (
  .P(P_2_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_2_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_9 (
  .P(P_2_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_2_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_2_10 (
  .P(P_2_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[50:34]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_0 (
  .P(P_3_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_1 (
  .P(P_3_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_2 (
  .P(P_3_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_3 (
  .P(P_3_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_4 (
  .P(P_3_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_5 (
  .P(P_3_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_6 (
  .P(P_3_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_7 (
  .P(P_3_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_8 (
  .P(P_3_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_3_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_9 (
  .P(P_3_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_3_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_3_10 (
  .P(P_3_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[67:51]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_0 (
  .P(P_4_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_1 (
  .P(P_4_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_2 (
  .P(P_4_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_3 (
  .P(P_4_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_4 (
  .P(P_4_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_5 (
  .P(P_4_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_6 (
  .P(P_4_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_7 (
  .P(P_4_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_8 (
  .P(P_4_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_4_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_9 (
  .P(P_4_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_4_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_4_10 (
  .P(P_4_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[84:68]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_0 (
  .P(P_5_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_1 (
  .P(P_5_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_2 (
  .P(P_5_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_3 (
  .P(P_5_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_4 (
  .P(P_5_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_5 (
  .P(P_5_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_6 (
  .P(P_5_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_7 (
  .P(P_5_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_8 (
  .P(P_5_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_5_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_9 (
  .P(P_5_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_5_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_5_10 (
  .P(P_5_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[101:85]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_0 (
  .P(P_6_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_1 (
  .P(P_6_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_2 (
  .P(P_6_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_3 (
  .P(P_6_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_4 (
  .P(P_6_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_5 (
  .P(P_6_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_6 (
  .P(P_6_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_7 (
  .P(P_6_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_8 (
  .P(P_6_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_6_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_9 (
  .P(P_6_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_6_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_6_10 (
  .P(P_6_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[118:102]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_0 (
  .P(P_7_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_1 (
  .P(P_7_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_2 (
  .P(P_7_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_3 (
  .P(P_7_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_4 (
  .P(P_7_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_5 (
  .P(P_7_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_6 (
  .P(P_7_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_7 (
  .P(P_7_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_8 (
  .P(P_7_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_7_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_9 (
  .P(P_7_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_7_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_7_10 (
  .P(P_7_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[135:119]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_0 (
  .P(P_8_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_1 (
  .P(P_8_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_2 (
  .P(P_8_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_3 (
  .P(P_8_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_4 (
  .P(P_8_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_5 (
  .P(P_8_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_6 (
  .P(P_8_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_7 (
  .P(P_8_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_8 (
  .P(P_8_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_8_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_9 (
  .P(P_8_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_8_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_8_10 (
  .P(P_8_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[152:136]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_0 (
  .P(P_9_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_1 (
  .P(P_9_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_2 (
  .P(P_9_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_3 (
  .P(P_9_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_4 (
  .P(P_9_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_5 (
  .P(P_9_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_6 (
  .P(P_9_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_7 (
  .P(P_9_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_8 (
  .P(P_9_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_9_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_9 (
  .P(P_9_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_9_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_9_10 (
  .P(P_9_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[169:153]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_0 (
  .P(P_10_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_1 (
  .P(P_10_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_2 (
  .P(P_10_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_3 (
  .P(P_10_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_4 (
  .P(P_10_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_5 (
  .P(P_10_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_6 (
  .P(P_10_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_7 (
  .P(P_10_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_8 (
  .P(P_10_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_10_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_9 (
  .P(P_10_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_10_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_10_10 (
  .P(P_10_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[186:170]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_0 (
  .P(P_11_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_1 (
  .P(P_11_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_2 (
  .P(P_11_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_3 (
  .P(P_11_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_4 (
  .P(P_11_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_5 (
  .P(P_11_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_6 (
  .P(P_11_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_7 (
  .P(P_11_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_8 (
  .P(P_11_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_11_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_9 (
  .P(P_11_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_11_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_11_10 (
  .P(P_11_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[203:187]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_0 (
  .P(P_12_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_1 (
  .P(P_12_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_2 (
  .P(P_12_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_3 (
  .P(P_12_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_4 (
  .P(P_12_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_5 (
  .P(P_12_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_6 (
  .P(P_12_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_7 (
  .P(P_12_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_8 (
  .P(P_12_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_12_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_9 (
  .P(P_12_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_12_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_12_10 (
  .P(P_12_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[220:204]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_0 (
  .P(P_13_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_1 (
  .P(P_13_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_2 (
  .P(P_13_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_3 (
  .P(P_13_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_4 (
  .P(P_13_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_5 (
  .P(P_13_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_6 (
  .P(P_13_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_7 (
  .P(P_13_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_8 (
  .P(P_13_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_13_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_9 (
  .P(P_13_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_13_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_13_10 (
  .P(P_13_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[237:221]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_0 (
  .P(P_14_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_1 (
  .P(P_14_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_2 (
  .P(P_14_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_3 (
  .P(P_14_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_4 (
  .P(P_14_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_5 (
  .P(P_14_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_6 (
  .P(P_14_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_7 (
  .P(P_14_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_8 (
  .P(P_14_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [42 : 0] P_14_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_9 (
  .P(P_14_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [34 : 0] P_14_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(18)        // Multiplier B-input bus width, 1-18
) MULT_14_10 (
  .P(P_14_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[254:238]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_0;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_0 (
  .P(P_15_0),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[23:0]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_1;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_1 (
  .P(P_15_1),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[47:24]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_2;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_2 (
  .P(P_15_2),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[71:48]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_3;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_3 (
  .P(P_15_3),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[95:72]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_4;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_4 (
  .P(P_15_4),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[119:96]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_5;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_5 (
  .P(P_15_5),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[143:120]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_6;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_6 (
  .P(P_15_6),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[167:144]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_7;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_7 (
  .P(P_15_7),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[191:168]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_8;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_8 (
  .P(P_15_8),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[215:192]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [26 : 0] P_15_9;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(25),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_9 (
  .P(P_15_9),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[239:216]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);

wire [18 : 0] P_15_10;

MULT #(
  .DEVICE("7SERIES"), // Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6","7SERIES"
  .LATENCY(3),        // Desired clock cycle latency, 0-4
  .WIDTH_A(17),       // Multiplier A-input bus width, 1-25
  .WIDTH_B(2)        // Multiplier B-input bus width, 1-18
) MULT_15_10 (
  .P(P_15_10),     // Multiplier output bus, width determined by WIDTH_P parameter
  .A({1'b0, mult_part_in0[255:240]}),     // Multiplier input A bus, width determined by WIDTH_A parameter
  .B({1'b0, mult_part_in1[255:255]}),     // Multiplier input B bus, width determined by WIDTH_B parameter
  .CE(CE),   // 1-bit active high input clock enable
  .CLK(clk), // 1-bit positive edge clock input
  .RST(rst)  // 1-bit input active high reset
);
always @(posedge clk)
    if (rst)
        begin
            mult_part_out00 <= 262'b0;
            mult_part_out01 <= 262'b0;
            mult_part_out02 <= 262'b0;
            mult_part_out03 <= 262'b0;
            mult_part_out04 <= 262'b0;
            mult_part_out05 <= 262'b0;
            mult_part_out06 <= 262'b0;
            mult_part_out07 <= 262'b0;
            mult_part_out08 <= 262'b0;
            mult_part_out09 <= 262'b0;
            mult_part_out10 <= 262'b0;
            mult_part_out11 <= 262'b0;
            mult_part_out12 <= 262'b0;
            mult_part_out13 <= 262'b0;
            mult_part_out14 <= 262'b0;
            mult_part_out15 <= 262'b0;
            mult_part_out16 <= 262'b0;
            mult_part_out17 <= 262'b0;
            mult_part_out18 <= 262'b0;
            mult_part_out19 <= 262'b0;
            mult_part_out20 <= 262'b0;
            mult_part_out21 <= 262'b0;
            mult_part_out22 <= 262'b0;
            mult_part_out23 <= 262'b0;
            mult_part_out24 <= 262'b0;
            mult_part_out25 <= 262'b0;
        end
    else
        begin
            mult_part_out00[0] <= P_0_0[0];
            mult_part_out00[1] <= P_0_0[1];
            mult_part_out00[2] <= P_0_0[2];
            mult_part_out00[3] <= P_0_0[3];
            mult_part_out00[4] <= P_0_0[4];
            mult_part_out00[5] <= P_0_0[5];
            mult_part_out00[6] <= P_0_0[6];
            mult_part_out00[7] <= P_0_0[7];
            mult_part_out00[8] <= P_0_0[8];
            mult_part_out00[9] <= P_0_0[9];
            mult_part_out00[10] <= P_0_0[10];
            mult_part_out00[11] <= P_0_0[11];
            mult_part_out00[12] <= P_0_0[12];
            mult_part_out00[13] <= P_0_0[13];
            mult_part_out00[14] <= P_0_0[14];
            mult_part_out00[15] <= P_0_0[15];
            mult_part_out00[16] <= P_0_0[16];
            mult_part_out00[17] <= P_1_0[0];
            mult_part_out00[18] <= P_1_0[1];
            mult_part_out00[19] <= P_0_0[19];
            mult_part_out00[20] <= P_1_0[3];
            mult_part_out00[21] <= P_0_0[21];
            mult_part_out00[22] <= P_1_0[5];
            mult_part_out00[23] <= P_0_0[23];
            mult_part_out00[24] <= P_1_0[7];
            mult_part_out00[25] <= P_0_0[25];
            mult_part_out00[26] <= P_0_0[26];
            mult_part_out00[27] <= P_0_1[3];
            mult_part_out00[28] <= P_0_0[28];
            mult_part_out00[29] <= P_0_0[29];
            mult_part_out00[30] <= P_0_1[6];
            mult_part_out00[31] <= P_1_0[14];
            mult_part_out00[32] <= P_0_0[32];
            mult_part_out00[33] <= P_1_0[16];
            mult_part_out00[34] <= P_2_0[0];
            mult_part_out00[35] <= P_2_0[1];
            mult_part_out00[36] <= P_1_0[19];
            mult_part_out00[37] <= P_1_0[20];
            mult_part_out00[38] <= P_0_0[38];
            mult_part_out00[39] <= P_1_0[22];
            mult_part_out00[40] <= P_0_1[16];
            mult_part_out00[41] <= P_1_1[0];
            mult_part_out00[42] <= P_1_1[1];
            mult_part_out00[43] <= P_1_1[2];
            mult_part_out00[44] <= P_2_0[10];
            mult_part_out00[45] <= P_1_0[28];
            mult_part_out00[46] <= P_2_0[12];
            mult_part_out00[47] <= P_1_0[30];
            mult_part_out00[48] <= P_1_1[7];
            mult_part_out00[49] <= P_1_0[32];
            mult_part_out00[50] <= P_1_1[9];
            mult_part_out00[51] <= P_1_0[34];
            mult_part_out00[52] <= P_0_2[4];
            mult_part_out00[53] <= P_3_0[2];
            mult_part_out00[54] <= P_1_0[37];
            mult_part_out00[55] <= P_3_0[4];
            mult_part_out00[56] <= P_2_0[22];
            mult_part_out00[57] <= P_2_0[23];
            mult_part_out00[58] <= P_0_2[10];
            mult_part_out00[59] <= P_2_0[25];
            mult_part_out00[60] <= P_0_2[12];
            mult_part_out00[61] <= P_1_1[20];
            mult_part_out00[62] <= P_2_0[28];
            mult_part_out00[63] <= P_0_2[15];
            mult_part_out00[64] <= P_0_1[40];
            mult_part_out00[65] <= P_3_0[14];
            mult_part_out00[66] <= P_3_0[15];
            mult_part_out00[67] <= P_3_0[16];
            mult_part_out00[68] <= P_1_1[27];
            mult_part_out00[69] <= P_2_1[11];
            mult_part_out00[70] <= P_4_0[2];
            mult_part_out00[71] <= P_0_2[23];
            mult_part_out00[72] <= P_1_1[31];
            mult_part_out00[73] <= P_3_0[22];
            mult_part_out00[74] <= P_0_3[2];
            mult_part_out00[75] <= P_1_1[34];
            mult_part_out00[76] <= P_4_0[8];
            mult_part_out00[77] <= P_1_2[12];
            mult_part_out00[78] <= P_0_2[30];
            mult_part_out00[79] <= P_1_1[38];
            mult_part_out00[80] <= P_0_3[8];
            mult_part_out00[81] <= P_3_0[30];
            mult_part_out00[82] <= P_2_2[0];
            mult_part_out00[83] <= P_2_2[1];
            mult_part_out00[84] <= P_0_2[36];
            mult_part_out00[85] <= P_0_2[37];
            mult_part_out00[86] <= P_2_1[28];
            mult_part_out00[87] <= P_1_2[22];
            mult_part_out00[88] <= P_0_2[40];
            mult_part_out00[89] <= P_2_2[7];
            mult_part_out00[90] <= P_2_2[8];
            mult_part_out00[91] <= P_0_3[19];
            mult_part_out00[92] <= P_5_0[7];
            mult_part_out00[93] <= P_2_1[35];
            mult_part_out00[94] <= P_2_1[36];
            mult_part_out00[95] <= P_4_0[27];
            mult_part_out00[96] <= P_2_1[38];
            mult_part_out00[97] <= P_2_1[39];
            mult_part_out00[98] <= P_2_1[40];
            mult_part_out00[99] <= P_4_0[31];
            mult_part_out00[100] <= P_4_0[32];
            mult_part_out00[101] <= P_5_0[16];
            mult_part_out00[102] <= P_4_0[34];
            mult_part_out00[103] <= P_6_0[1];
            mult_part_out00[104] <= P_0_3[32];
            mult_part_out00[105] <= P_0_3[33];
            mult_part_out00[106] <= P_2_3[0];
            mult_part_out00[107] <= P_2_3[1];
            mult_part_out00[108] <= P_3_1[33];
            mult_part_out00[109] <= P_4_1[17];
            mult_part_out00[110] <= P_2_3[4];
            mult_part_out00[111] <= P_5_0[26];
            mult_part_out00[112] <= P_2_2[30];
            mult_part_out00[113] <= P_2_3[7];
            mult_part_out00[114] <= P_1_4[1];
            mult_part_out00[115] <= P_3_1[40];
            mult_part_out00[116] <= P_1_4[3];
            mult_part_out00[117] <= P_5_1[8];
            mult_part_out00[118] <= P_2_3[12];
            mult_part_out00[119] <= P_5_0[34];
            mult_part_out00[120] <= P_1_3[31];
            mult_part_out00[121] <= P_7_0[2];
            mult_part_out00[122] <= P_5_1[13];
            mult_part_out00[123] <= P_5_0[38];
            mult_part_out00[124] <= P_5_0[39];
            mult_part_out00[125] <= P_4_2[9];
            mult_part_out00[126] <= P_3_2[27];
            mult_part_out00[127] <= P_4_1[35];
            mult_part_out00[128] <= P_5_1[19];
            mult_part_out00[129] <= P_5_1[20];
            mult_part_out00[130] <= P_0_4[34];
            mult_part_out00[131] <= P_0_4[35];
            mult_part_out00[132] <= P_6_1[6];
            mult_part_out00[133] <= P_6_0[31];
            mult_part_out00[134] <= P_5_2[1];
            mult_part_out00[135] <= P_3_2[36];
            mult_part_out00[136] <= P_1_4[23];
            mult_part_out00[137] <= P_5_1[28];
            mult_part_out00[138] <= P_1_5[1];
            mult_part_out00[139] <= P_7_0[20];
            mult_part_out00[140] <= P_5_2[7];
            mult_part_out00[141] <= P_7_0[22];
            mult_part_out00[142] <= P_6_0[40];
            mult_part_out00[143] <= P_4_3[3];
            mult_part_out00[144] <= P_1_4[31];
            mult_part_out00[145] <= P_7_0[26];
            mult_part_out00[146] <= P_1_4[33];
            mult_part_out00[147] <= P_5_1[38];
            mult_part_out00[148] <= P_7_1[5];
            mult_part_out00[149] <= P_1_5[12];
            mult_part_out00[150] <= P_7_0[31];
            mult_part_out00[151] <= P_1_5[14];
            mult_part_out00[152] <= P_0_5[32];
            mult_part_out00[153] <= P_0_5[33];
            mult_part_out00[154] <= P_5_2[21];
            mult_part_out00[155] <= P_0_6[11];
            mult_part_out00[156] <= P_6_1[30];
            mult_part_out00[157] <= P_9_0[4];
            mult_part_out00[158] <= P_5_2[25];
            mult_part_out00[159] <= P_7_0[40];
            mult_part_out00[160] <= P_6_1[34];
            mult_part_out00[161] <= P_7_1[18];
            mult_part_out00[162] <= P_2_4[32];
            mult_part_out00[163] <= P_2_4[33];
            mult_part_out00[164] <= P_8_1[4];
            mult_part_out00[165] <= P_2_4[35];
            mult_part_out00[166] <= P_2_5[12];
            mult_part_out00[167] <= P_6_2[17];
            mult_part_out00[168] <= P_8_1[8];
            mult_part_out00[169] <= P_2_4[39];
            mult_part_out00[170] <= P_6_2[20];
            mult_part_out00[171] <= P_6_2[21];
            mult_part_out00[172] <= P_0_7[4];
            mult_part_out00[173] <= P_8_1[13];
            mult_part_out00[174] <= P_7_1[31];
            mult_part_out00[175] <= P_7_2[8];
            mult_part_out00[176] <= P_0_7[8];
            mult_part_out00[177] <= P_3_5[6];
            mult_part_out00[178] <= P_6_3[4];
            mult_part_out00[179] <= P_6_3[5];
            mult_part_out00[180] <= P_2_6[2];
            mult_part_out00[181] <= P_0_6[37];
            mult_part_out00[182] <= P_2_6[4];
            mult_part_out00[183] <= P_9_1[6];
            mult_part_out00[184] <= P_8_2[0];
            mult_part_out00[185] <= P_8_1[25];
            mult_part_out00[186] <= P_8_1[26];
            mult_part_out00[187] <= P_9_0[34];
            mult_part_out00[188] <= P_5_3[31];
            mult_part_out00[189] <= P_5_3[32];
            mult_part_out00[190] <= P_3_5[19];
            mult_part_out00[191] <= P_6_3[17];
            mult_part_out00[192] <= P_5_3[35];
            mult_part_out00[193] <= P_2_6[15];
            mult_part_out00[194] <= P_7_2[27];
            mult_part_out00[195] <= P_1_7[10];
            mult_part_out00[196] <= P_6_3[22];
            mult_part_out00[197] <= P_4_4[33];
            mult_part_out00[198] <= P_10_1[4];
            mult_part_out00[199] <= P_2_6[21];
            mult_part_out00[200] <= P_10_1[6];
            mult_part_out00[201] <= P_3_6[6];
            mult_part_out00[202] <= P_8_2[18];
            mult_part_out00[203] <= P_7_2[36];
            mult_part_out00[204] <= P_11_0[17];
            mult_part_out00[205] <= P_0_8[13];
            mult_part_out00[206] <= P_0_7[38];
            mult_part_out00[207] <= P_11_0[20];
            mult_part_out00[208] <= P_10_0[38];
            mult_part_out00[209] <= P_0_8[17];
            mult_part_out00[210] <= P_0_8[18];
            mult_part_out00[211] <= P_7_3[20];
            mult_part_out00[212] <= P_0_8[20];
            mult_part_out00[213] <= P_5_5[8];
            mult_part_out00[214] <= P_5_4[33];
            mult_part_out00[215] <= P_11_0[28];
            mult_part_out00[216] <= P_3_6[21];
            mult_part_out00[217] <= P_0_8[25];
            mult_part_out00[218] <= P_11_1[7];
            mult_part_out00[219] <= P_4_6[7];
            mult_part_out00[220] <= P_1_8[11];
            mult_part_out00[221] <= P_3_6[26];
            mult_part_out00[222] <= P_4_6[10];
            mult_part_out00[223] <= P_3_7[4];
            mult_part_out00[224] <= P_12_0[20];
            mult_part_out00[225] <= P_13_0[4];
            mult_part_out00[226] <= P_2_8[0];
            mult_part_out00[227] <= P_10_2[9];
            mult_part_out00[228] <= P_12_1[0];
            mult_part_out00[229] <= P_11_1[18];
            mult_part_out00[230] <= P_3_6[35];
            mult_part_out00[231] <= P_10_1[37];
            mult_part_out00[232] <= P_6_5[10];
            mult_part_out00[233] <= P_12_1[5];
            mult_part_out00[234] <= P_13_0[13];
            mult_part_out00[235] <= P_11_2[0];
            mult_part_out00[236] <= P_9_3[11];
            mult_part_out00[237] <= P_12_1[9];
            mult_part_out00[238] <= P_13_0[17];
            mult_part_out00[239] <= P_8_3[31];
            mult_part_out00[240] <= P_11_2[5];
            mult_part_out00[241] <= P_11_2[6];
            mult_part_out00[242] <= P_0_9[26];
            mult_part_out00[243] <= P_8_3[35];
            mult_part_out00[244] <= P_3_8[1];
            mult_part_out00[245] <= P_10_3[3];
            mult_part_out00[246] <= P_7_5[7];
            mult_part_out00[247] <= P_9_3[22];
            mult_part_out00[248] <= P_9_3[23];
            mult_part_out00[249] <= P_6_6[3];
            mult_part_out00[250] <= P_11_1[39];
            mult_part_out00[251] <= P_7_4[36];
            mult_part_out00[252] <= P_12_1[24];
            mult_part_out00[253] <= P_3_7[34];
            mult_part_out00[254] <= P_4_7[18];
            mult_part_out00[255] <= P_2_9[5];
            mult_part_out00[256] <= P_10_3[14];
            mult_part_out00[257] <= P_1_9[24];
            mult_part_out00[258] <= P_5_7[5];
            mult_part_out00[259] <= P_9_3[34];
            mult_part_out00[260] <= P_13_0[39];
            mult_part_out00[261] <= P_7_5[22];
            mult_part_out00[262] <= P_15_0[7];
            mult_part_out00[263] <= P_1_9[30];
            mult_part_out00[264] <= P_1_10[7];
            mult_part_out00[265] <= P_9_4[16];
            mult_part_out00[266] <= P_12_2[14];
            mult_part_out00[267] <= P_4_8[7];
            mult_part_out00[268] <= P_1_9[35];
            mult_part_out00[269] <= P_10_4[3];
            mult_part_out00[270] <= P_10_3[28];
            mult_part_out00[271] <= P_1_10[14];
            mult_part_out00[272] <= P_5_7[19];
            mult_part_out00[273] <= P_2_9[23];
            mult_part_out00[274] <= P_8_5[18];
            mult_part_out00[275] <= P_2_10[1];
            mult_part_out00[276] <= P_9_5[3];
            mult_part_out00[277] <= P_3_8[34];
            mult_part_out00[278] <= P_6_6[32];
            mult_part_out00[279] <= P_13_1[34];
            mult_part_out00[280] <= P_4_8[20];
            mult_part_out00[281] <= P_5_7[28];
            mult_part_out00[282] <= P_11_3[23];
            mult_part_out00[283] <= P_3_8[40];
            mult_part_out00[284] <= P_10_4[18];
            mult_part_out00[285] <= P_3_9[18];
            mult_part_out00[286] <= P_14_2[0];
            mult_part_out00[287] <= P_1_10[30];
            mult_part_out00[288] <= P_7_6[25];
            mult_part_out00[289] <= P_11_3[30];
            mult_part_out00[290] <= P_10_4[24];
            mult_part_out00[291] <= P_10_5[1];
            mult_part_out00[292] <= P_12_2[40];
            mult_part_out00[293] <= P_10_4[27];
            mult_part_out00[294] <= P_9_5[21];
            mult_part_out00[295] <= P_13_2[26];
            mult_part_out00[296] <= P_6_7[26];
            mult_part_out00[297] <= P_3_9[30];
            mult_part_out00[298] <= P_4_8[38];
            mult_part_out00[299] <= P_7_7[12];
            mult_part_out00[300] <= P_9_6[3];
            mult_part_out00[301] <= P_15_1[22];
            mult_part_out00[302] <= P_9_5[29];
            mult_part_out00[303] <= P_3_9[36];
            mult_part_out00[304] <= P_8_6[24];
            mult_part_out00[305] <= P_6_7[35];
            mult_part_out00[306] <= P_8_6[26];
            mult_part_out00[307] <= P_13_3[14];
            mult_part_out00[308] <= P_6_7[38];
            mult_part_out00[309] <= P_3_10[18];
            mult_part_out00[310] <= P_14_3[0];
            mult_part_out00[311] <= P_3_10[20];
            mult_part_out00[312] <= P_12_4[12];
            mult_part_out00[313] <= P_7_7[26];
            mult_part_out00[314] <= P_9_6[17];
            mult_part_out00[315] <= P_6_8[21];
            mult_part_out00[316] <= P_5_9[15];
            mult_part_out00[317] <= P_15_2[14];
            mult_part_out00[318] <= P_13_3[25];
            mult_part_out00[319] <= P_11_4[36];
            mult_part_out00[320] <= P_9_6[23];
            mult_part_out00[321] <= P_13_3[28];
            mult_part_out00[322] <= P_7_8[11];
            mult_part_out00[323] <= P_10_6[9];
            mult_part_out00[324] <= P_7_8[13];
            mult_part_out00[325] <= P_7_8[14];
            mult_part_out00[326] <= P_14_2[40];
            mult_part_out00[327] <= P_12_5[3];
            mult_part_out00[328] <= P_14_3[18];
            mult_part_out00[329] <= P_5_10[4];
            mult_part_out00[330] <= P_4_10[22];
            mult_part_out00[331] <= P_13_4[14];
            mult_part_out00[332] <= P_11_5[25];
            mult_part_out00[333] <= P_10_6[19];
            mult_part_out00[334] <= P_14_4[0];
            mult_part_out00[335] <= P_8_7[31];
            mult_part_out00[336] <= P_9_6[39];
            mult_part_out00[337] <= P_10_6[23];
            mult_part_out00[338] <= P_12_4[38];
            mult_part_out00[339] <= P_8_7[35];
            mult_part_out00[340] <= P_15_3[13];
            mult_part_out00[341] <= P_13_4[24];
            mult_part_out00[342] <= P_15_3[15];
            mult_part_out00[343] <= P_13_4[26];
            mult_part_out00[344] <= P_11_5[37];
            mult_part_out00[345] <= P_7_8[34];
            mult_part_out00[346] <= P_6_10[4];
            mult_part_out00[347] <= P_10_6[33];
            mult_part_out00[348] <= P_14_3[38];
            mult_part_out00[349] <= P_6_10[7];
            mult_part_out00[350] <= P_15_3[23];
            mult_part_out00[351] <= P_12_6[3];
            mult_part_out00[352] <= P_15_4[1];
            mult_part_out00[353] <= P_5_10[28];
            mult_part_out00[354] <= P_6_9[36];
            mult_part_out00[355] <= P_11_7[0];
            mult_part_out00[356] <= P_5_10[31];
            mult_part_out00[357] <= P_14_4[23];
            mult_part_out00[358] <= P_12_6[10];
            mult_part_out00[359] <= P_7_10[0];
            mult_part_out00[360] <= P_10_7[22];
            mult_part_out00[361] <= P_15_4[10];
            mult_part_out00[362] <= P_10_8[0];
            mult_part_out00[363] <= P_10_7[25];
            mult_part_out00[364] <= P_8_8[36];
            mult_part_out00[365] <= P_8_8[37];
            mult_part_out00[366] <= P_14_5[8];
            mult_part_out00[367] <= P_11_6[36];
            mult_part_out00[368] <= P_14_5[10];
            mult_part_out00[369] <= P_9_8[24];
            mult_part_out00[370] <= P_6_10[28];
            mult_part_out00[371] <= P_9_8[26];
            mult_part_out00[372] <= P_11_7[17];
            mult_part_out00[373] <= P_12_7[1];
            mult_part_out00[374] <= P_10_7[36];
            mult_part_out00[375] <= P_10_7[37];
            mult_part_out00[376] <= P_13_6[11];
            mult_part_out00[377] <= P_15_5[2];
            mult_part_out00[378] <= P_14_5[20];
            mult_part_out00[379] <= P_13_6[14];
            mult_part_out00[380] <= P_8_9[28];
            mult_part_out00[381] <= P_11_7[26];
            mult_part_out00[382] <= P_12_7[10];
            mult_part_out00[383] <= P_11_7[28];
            mult_part_out00[384] <= P_15_5[9];
            mult_part_out00[385] <= P_8_9[33];
            mult_part_out00[386] <= P_13_6[21];
            mult_part_out00[387] <= P_14_6[5];
            mult_part_out00[388] <= P_10_9[2];
            mult_part_out00[389] <= P_8_10[13];
            mult_part_out00[390] <= P_10_9[4];
            mult_part_out00[391] <= P_8_9[39];
            mult_part_out00[392] <= P_8_9[40];
            mult_part_out00[393] <= P_15_5[18];
            mult_part_out00[394] <= P_8_10[18];
            mult_part_out00[395] <= P_11_7[40];
            mult_part_out00[396] <= P_12_8[0];
            mult_part_out00[397] <= P_12_7[25];
            mult_part_out00[398] <= P_14_6[16];
            mult_part_out00[399] <= P_12_8[3];
            mult_part_out00[400] <= P_11_8[21];
            mult_part_out00[401] <= P_15_6[2];
            mult_part_out00[402] <= P_13_6[37];
            mult_part_out00[403] <= P_9_9[34];
            mult_part_out00[404] <= P_12_7[32];
            mult_part_out00[405] <= P_10_9[19];
            mult_part_out00[406] <= P_15_6[7];
            mult_part_out00[407] <= P_15_6[8];
            mult_part_out00[408] <= P_12_7[36];
            mult_part_out00[409] <= P_14_7[3];
            mult_part_out00[410] <= P_11_9[7];
            mult_part_out00[411] <= P_10_9[25];
            mult_part_out00[412] <= P_11_9[9];
            mult_part_out00[413] <= P_9_10[20];
            mult_part_out00[414] <= P_14_6[32];
            mult_part_out00[415] <= P_11_9[12];
            mult_part_out00[416] <= P_9_10[23];
            mult_part_out00[417] <= P_15_6[18];
            mult_part_out00[418] <= P_12_8[22];
            mult_part_out00[419] <= P_11_8[40];
            mult_part_out00[420] <= P_14_6[38];
            mult_part_out00[421] <= P_14_6[39];
            mult_part_out00[422] <= P_14_7[16];
            mult_part_out00[423] <= P_14_7[17];
            mult_part_out00[424] <= P_12_9[4];
            mult_part_out00[425] <= P_10_10[15];
            mult_part_out00[426] <= P_10_9[40];
            mult_part_out00[427] <= P_11_9[24];
            mult_part_out00[428] <= P_10_10[18];
            mult_part_out00[429] <= P_10_10[19];
            mult_part_out00[430] <= P_15_7[7];
            mult_part_out00[431] <= P_11_9[28];
            mult_part_out00[432] <= P_11_10[5];
            mult_part_out00[433] <= P_10_10[23];
            mult_part_out00[434] <= P_12_8[38];
            mult_part_out00[435] <= P_12_9[15];
            mult_part_out00[436] <= P_11_9[33];
            mult_part_out00[437] <= P_13_8[24];
            mult_part_out00[438] <= P_14_8[8];
            mult_part_out00[439] <= P_14_8[9];
            mult_part_out00[440] <= P_11_9[37];
            mult_part_out00[441] <= P_13_8[28];
            mult_part_out00[442] <= P_10_10[32];
            mult_part_out00[443] <= P_11_10[16];
            mult_part_out00[444] <= P_11_10[17];
            mult_part_out00[445] <= P_13_9[8];
            mult_part_out00[446] <= P_15_7[23];
            mult_part_out00[447] <= P_14_8[17];
            mult_part_out00[448] <= P_14_8[18];
            mult_part_out00[449] <= P_15_8[2];
            mult_part_out00[450] <= P_13_8[37];
            mult_part_out00[451] <= P_14_8[21];
            mult_part_out00[452] <= P_11_10[25];
            mult_part_out00[453] <= P_11_10[26];
            mult_part_out00[454] <= P_15_8[7];
            mult_part_out00[455] <= P_14_8[25];
            mult_part_out00[456] <= P_14_9[2];
            mult_part_out00[457] <= P_15_8[10];
            mult_part_out00[458] <= P_13_9[21];
            mult_part_out00[459] <= P_12_10[15];
            mult_part_out00[460] <= P_12_10[16];
            mult_part_out00[461] <= P_14_8[31];
            mult_part_out00[462] <= P_12_10[18];
            mult_part_out00[463] <= P_14_9[9];
            mult_part_out00[464] <= P_15_8[17];
            mult_part_out00[465] <= P_14_8[35];
            mult_part_out00[466] <= P_15_8[19];
            mult_part_out00[467] <= P_15_8[20];
            mult_part_out00[468] <= P_13_10[7];
            mult_part_out00[469] <= P_14_8[39];
            mult_part_out00[470] <= P_13_10[9];
            mult_part_out00[471] <= P_12_10[27];
            mult_part_out00[472] <= P_14_9[18];
            mult_part_out00[473] <= P_12_10[29];
            mult_part_out00[474] <= P_13_10[13];
            mult_part_out00[475] <= P_12_10[31];
            mult_part_out00[476] <= P_13_10[15];
            mult_part_out00[477] <= P_13_9[40];
            mult_part_out00[478] <= P_14_10[0];
            mult_part_out00[479] <= P_14_10[1];
            mult_part_out00[480] <= P_14_9[26];
            mult_part_out00[481] <= P_14_9[27];
            mult_part_out00[482] <= P_15_9[11];
            mult_part_out00[483] <= P_14_9[29];
            mult_part_out00[484] <= P_14_10[6];
            mult_part_out00[485] <= P_15_9[14];
            mult_part_out00[486] <= P_13_10[25];
            mult_part_out00[487] <= P_13_10[26];
            mult_part_out00[488] <= P_15_9[17];
            mult_part_out00[489] <= P_14_10[11];
            mult_part_out00[490] <= P_14_10[12];
            mult_part_out00[491] <= P_14_9[37];
            mult_part_out00[492] <= P_14_10[14];
            mult_part_out00[493] <= P_14_10[15];
            mult_part_out00[494] <= P_15_9[23];
            mult_part_out00[495] <= P_15_10[0];
            mult_part_out00[496] <= P_15_10[1];
            mult_part_out00[497] <= P_14_10[19];
            mult_part_out00[498] <= P_15_10[3];
            mult_part_out00[499] <= P_14_10[21];
            mult_part_out00[500] <= P_15_10[5];
            mult_part_out00[501] <= P_14_10[23];
            mult_part_out00[502] <= P_15_10[7];
            mult_part_out00[503] <= P_14_10[25];
            mult_part_out00[504] <= P_14_10[26];
            mult_part_out00[505] <= P_14_10[27];
            mult_part_out00[506] <= P_15_10[11];
            mult_part_out00[507] <= P_14_10[29];
            mult_part_out00[508] <= P_15_10[13];
            mult_part_out00[509] <= P_14_10[31];
            mult_part_out00[510] <= P_14_10[32];
            mult_part_out00[511] <= P_15_10[16];

            mult_part_out01[17] <= P_0_0[17];
            mult_part_out01[18] <= P_0_0[18];
            mult_part_out01[19] <= P_1_0[2];
            mult_part_out01[20] <= P_0_0[20];
            mult_part_out01[21] <= P_1_0[4];
            mult_part_out01[22] <= P_0_0[22];
            mult_part_out01[23] <= P_1_0[6];
            mult_part_out01[24] <= P_0_0[24];
            mult_part_out01[25] <= P_0_1[1];
            mult_part_out01[26] <= P_0_1[2];
            mult_part_out01[27] <= P_1_0[10];
            mult_part_out01[28] <= P_0_1[4];
            mult_part_out01[29] <= P_0_1[5];
            mult_part_out01[30] <= P_1_0[13];
            mult_part_out01[31] <= P_0_0[31];
            mult_part_out01[32] <= P_0_1[8];
            mult_part_out01[33] <= P_0_0[33];
            mult_part_out01[34] <= P_0_0[34];
            mult_part_out01[35] <= P_0_0[35];
            mult_part_out01[36] <= P_2_0[2];
            mult_part_out01[37] <= P_2_0[3];
            mult_part_out01[38] <= P_0_1[14];
            mult_part_out01[39] <= P_2_0[5];
            mult_part_out01[40] <= P_1_0[23];
            mult_part_out01[41] <= P_0_1[17];
            mult_part_out01[42] <= P_1_0[25];
            mult_part_out01[43] <= P_0_1[19];
            mult_part_out01[44] <= P_0_1[20];
            mult_part_out01[45] <= P_0_1[21];
            mult_part_out01[46] <= P_0_1[22];
            mult_part_out01[47] <= P_0_1[23];
            mult_part_out01[48] <= P_0_2[0];
            mult_part_out01[49] <= P_0_2[1];
            mult_part_out01[50] <= P_2_0[16];
            mult_part_out01[51] <= P_1_1[10];
            mult_part_out01[52] <= P_1_0[35];
            mult_part_out01[53] <= P_0_1[29];
            mult_part_out01[54] <= P_0_2[6];
            mult_part_out01[55] <= P_1_1[14];
            mult_part_out01[56] <= P_0_2[8];
            mult_part_out01[57] <= P_3_0[6];
            mult_part_out01[58] <= P_3_0[7];
            mult_part_out01[59] <= P_0_2[11];
            mult_part_out01[60] <= P_2_0[26];
            mult_part_out01[61] <= P_2_1[3];
            mult_part_out01[62] <= P_0_1[38];
            mult_part_out01[63] <= P_0_1[39];
            mult_part_out01[64] <= P_3_0[13];
            mult_part_out01[65] <= P_2_1[7];
            mult_part_out01[66] <= P_1_1[25];
            mult_part_out01[67] <= P_2_0[33];
            mult_part_out01[68] <= P_1_2[3];
            mult_part_out01[69] <= P_0_2[21];
            mult_part_out01[70] <= P_2_1[12];
            mult_part_out01[71] <= P_1_1[30];
            mult_part_out01[72] <= P_2_0[38];
            mult_part_out01[73] <= P_2_0[39];
            mult_part_out01[74] <= P_1_1[33];
            mult_part_out01[75] <= P_3_1[0];
            mult_part_out01[76] <= P_1_1[35];
            mult_part_out01[77] <= P_2_1[19];
            mult_part_out01[78] <= P_2_1[20];
            mult_part_out01[79] <= P_0_2[31];
            mult_part_out01[80] <= P_3_0[29];
            mult_part_out01[81] <= P_0_2[33];
            mult_part_out01[82] <= P_4_0[14];
            mult_part_out01[83] <= P_3_0[32];
            mult_part_out01[84] <= P_0_3[12];
            mult_part_out01[85] <= P_5_0[0];
            mult_part_out01[86] <= P_0_3[14];
            mult_part_out01[87] <= P_5_0[2];
            mult_part_out01[88] <= P_3_0[37];
            mult_part_out01[89] <= P_4_0[21];
            mult_part_out01[90] <= P_4_0[22];
            mult_part_out01[91] <= P_3_0[40];
            mult_part_out01[92] <= P_4_0[24];
            mult_part_out01[93] <= P_2_2[11];
            mult_part_out01[94] <= P_5_0[9];
            mult_part_out01[95] <= P_1_3[6];
            mult_part_out01[96] <= P_4_0[28];
            mult_part_out01[97] <= P_4_0[29];
            mult_part_out01[98] <= P_1_2[33];
            mult_part_out01[99] <= P_2_2[17];
            mult_part_out01[100] <= P_3_1[25];
            mult_part_out01[101] <= P_4_1[9];
            mult_part_out01[102] <= P_3_1[27];
            mult_part_out01[103] <= P_3_2[4];
            mult_part_out01[104] <= P_4_1[12];
            mult_part_out01[105] <= P_1_3[16];
            mult_part_out01[106] <= P_5_0[21];
            mult_part_out01[107] <= P_6_0[5];
            mult_part_out01[108] <= P_6_0[6];
            mult_part_out01[109] <= P_2_3[3];
            mult_part_out01[110] <= P_3_2[11];
            mult_part_out01[111] <= P_3_1[36];
            mult_part_out01[112] <= P_3_2[13];
            mult_part_out01[113] <= P_2_2[31];
            mult_part_out01[114] <= P_0_4[18];
            mult_part_out01[115] <= P_0_4[19];
            mult_part_out01[116] <= P_1_3[27];
            mult_part_out01[117] <= P_4_1[25];
            mult_part_out01[118] <= P_3_2[19];
            mult_part_out01[119] <= P_1_3[30];
            mult_part_out01[120] <= P_2_3[14];
            mult_part_out01[121] <= P_0_4[25];
            mult_part_out01[122] <= P_7_0[3];
            mult_part_out01[123] <= P_4_1[31];
            mult_part_out01[124] <= P_0_4[28];
            mult_part_out01[125] <= P_6_0[23];
            mult_part_out01[126] <= P_0_5[6];
            mult_part_out01[127] <= P_5_1[18];
            mult_part_out01[128] <= P_4_1[36];
            mult_part_out01[129] <= P_0_5[9];
            mult_part_out01[130] <= P_0_5[10];
            mult_part_out01[131] <= P_7_0[12];
            mult_part_out01[132] <= P_2_4[2];
            mult_part_out01[133] <= P_1_4[20];
            mult_part_out01[134] <= P_1_4[21];
            mult_part_out01[135] <= P_7_0[16];
            mult_part_out01[136] <= P_5_2[3];
            mult_part_out01[137] <= P_1_5[0];
            mult_part_out01[138] <= P_2_3[32];
            mult_part_out01[139] <= P_2_4[9];
            mult_part_out01[140] <= P_6_1[14];
            mult_part_out01[141] <= P_8_0[5];
            mult_part_out01[142] <= P_5_2[9];
            mult_part_out01[143] <= P_4_2[27];
            mult_part_out01[144] <= P_3_3[21];
            mult_part_out01[145] <= P_1_4[32];
            mult_part_out01[146] <= P_3_3[23];
            mult_part_out01[147] <= P_8_0[11];
            mult_part_out01[148] <= P_4_2[32];
            mult_part_out01[149] <= P_5_2[16];
            mult_part_out01[150] <= P_2_4[20];
            mult_part_out01[151] <= P_6_2[1];
            mult_part_out01[152] <= P_6_2[2];
            mult_part_out01[153] <= P_0_6[9];
            mult_part_out01[154] <= P_4_2[38];
            mult_part_out01[155] <= P_5_2[22];
            mult_part_out01[156] <= P_0_5[36];
            mult_part_out01[157] <= P_4_3[17];
            mult_part_out01[158] <= P_5_3[1];
            mult_part_out01[159] <= P_7_1[16];
            mult_part_out01[160] <= P_9_0[7];
            mult_part_out01[161] <= P_6_1[35];
            mult_part_out01[162] <= P_1_6[1];
            mult_part_out01[163] <= P_1_5[26];
            mult_part_out01[164] <= P_5_3[7];
            mult_part_out01[165] <= P_3_4[18];
            mult_part_out01[166] <= P_8_1[6];
            mult_part_out01[167] <= P_9_0[14];
            mult_part_out01[168] <= P_1_5[31];
            mult_part_out01[169] <= P_9_0[16];
            mult_part_out01[170] <= P_2_4[40];
            mult_part_out01[171] <= P_4_4[7];
            mult_part_out01[172] <= P_7_2[5];
            mult_part_out01[173] <= P_9_0[20];
            mult_part_out01[174] <= P_6_3[0];
            mult_part_out01[175] <= P_10_0[5];
            mult_part_out01[176] <= P_8_1[16];
            mult_part_out01[177] <= P_9_1[0];
            mult_part_out01[178] <= P_5_3[21];
            mult_part_out01[179] <= P_4_4[15];
            mult_part_out01[180] <= P_10_0[10];
            mult_part_out01[181] <= P_1_6[20];
            mult_part_out01[182] <= P_4_4[18];
            mult_part_out01[183] <= P_3_5[12];
            mult_part_out01[184] <= P_1_6[23];
            mult_part_out01[185] <= P_8_2[1];
            mult_part_out01[186] <= P_10_0[16];
            mult_part_out01[187] <= P_3_4[40];
            mult_part_out01[188] <= P_6_2[38];
            mult_part_out01[189] <= P_6_3[15];
            mult_part_out01[190] <= P_1_6[29];
            mult_part_out01[191] <= P_9_1[14];
            mult_part_out01[192] <= P_7_2[25];
            mult_part_out01[193] <= P_5_3[36];
            mult_part_out01[194] <= P_9_1[17];
            mult_part_out01[195] <= P_7_3[4];
            mult_part_out01[196] <= P_5_3[39];
            mult_part_out01[197] <= P_5_3[40];
            mult_part_out01[198] <= P_7_3[7];
            mult_part_out01[199] <= P_9_1[22];
            mult_part_out01[200] <= P_4_4[36];
            mult_part_out01[201] <= P_4_4[37];
            mult_part_out01[202] <= P_9_2[1];
            mult_part_out01[203] <= P_9_1[26];
            mult_part_out01[204] <= P_9_2[3];
            mult_part_out01[205] <= P_10_0[35];
            mult_part_out01[206] <= P_1_7[21];
            mult_part_out01[207] <= P_6_4[9];
            mult_part_out01[208] <= P_4_5[20];
            mult_part_out01[209] <= P_1_8[0];
            mult_part_out01[210] <= P_2_7[8];
            mult_part_out01[211] <= P_0_8[19];
            mult_part_out01[212] <= P_6_4[14];
            mult_part_out01[213] <= P_11_0[26];
            mult_part_out01[214] <= P_1_7[29];
            mult_part_out01[215] <= P_8_2[31];
            mult_part_out01[216] <= P_4_6[4];
            mult_part_out01[217] <= P_7_4[2];
            mult_part_out01[218] <= P_2_7[16];
            mult_part_out01[219] <= P_7_4[4];
            mult_part_out01[220] <= P_11_1[9];
            mult_part_out01[221] <= P_10_1[27];
            mult_part_out01[222] <= P_9_2[21];
            mult_part_out01[223] <= P_8_3[15];
            mult_part_out01[224] <= P_8_3[16];
            mult_part_out01[225] <= P_0_9[9];
            mult_part_out01[226] <= P_2_7[24];
            mult_part_out01[227] <= P_4_6[15];
            mult_part_out01[228] <= P_3_7[9];
            mult_part_out01[229] <= P_4_6[17];
            mult_part_out01[230] <= P_12_1[2];
            mult_part_out01[231] <= P_0_9[15];
            mult_part_out01[232] <= P_6_4[34];
            mult_part_out01[233] <= P_4_6[21];
            mult_part_out01[234] <= P_10_1[40];
            mult_part_out01[235] <= P_9_3[10];
            mult_part_out01[236] <= P_7_4[21];
            mult_part_out01[237] <= P_11_2[2];
            mult_part_out01[238] <= P_10_2[20];
            mult_part_out01[239] <= P_11_1[28];
            mult_part_out01[240] <= P_8_3[32];
            mult_part_out01[241] <= P_11_1[30];
            mult_part_out01[242] <= P_12_1[14];
            mult_part_out01[243] <= P_12_1[15];
            mult_part_out01[244] <= P_0_9[28];
            mult_part_out01[245] <= P_14_0[7];
            mult_part_out01[246] <= P_0_9[30];
            mult_part_out01[247] <= P_0_10[7];
            mult_part_out01[248] <= P_11_1[37];
            mult_part_out01[249] <= P_8_4[17];
            mult_part_out01[250] <= P_3_8[7];
            mult_part_out01[251] <= P_7_5[12];
            mult_part_out01[252] <= P_13_1[7];
            mult_part_out01[253] <= P_12_2[1];
            mult_part_out01[254] <= P_8_4[22];
            mult_part_out01[255] <= P_6_5[33];
            mult_part_out01[256] <= P_6_6[10];
            mult_part_out01[257] <= P_9_3[32];
            mult_part_out01[258] <= P_0_10[18];
            mult_part_out01[259] <= P_1_10[2];
            mult_part_out01[260] <= P_9_4[11];
            mult_part_out01[261] <= P_6_5[39];
            mult_part_out01[262] <= P_4_8[2];
            mult_part_out01[263] <= P_14_1[1];
            mult_part_out01[264] <= P_14_1[2];
            mult_part_out01[265] <= P_1_9[32];
            mult_part_out01[266] <= P_6_6[20];
            mult_part_out01[267] <= P_4_7[31];
            mult_part_out01[268] <= P_0_10[28];
            mult_part_out01[269] <= P_13_2[0];
            mult_part_out01[270] <= P_11_3[11];
            mult_part_out01[271] <= P_10_3[29];
            mult_part_out01[272] <= P_4_8[12];
            mult_part_out01[273] <= P_4_7[37];
            mult_part_out01[274] <= P_1_10[17];
            mult_part_out01[275] <= P_13_1[30];
            mult_part_out01[276] <= P_11_3[17];
            mult_part_out01[277] <= P_4_8[17];
            mult_part_out01[278] <= P_12_3[2];
            mult_part_out01[279] <= P_8_5[23];
            mult_part_out01[280] <= P_3_8[37];
            mult_part_out01[281] <= P_8_5[25];
            mult_part_out01[282] <= P_2_9[32];
            mult_part_out01[283] <= P_6_6[37];
            mult_part_out01[284] <= P_9_4[35];
            mult_part_out01[285] <= P_7_6[22];
            mult_part_out01[286] <= P_9_4[37];
            mult_part_out01[287] <= P_7_7[0];
            mult_part_out01[288] <= P_14_1[26];
            mult_part_out01[289] <= P_13_2[20];
            mult_part_out01[290] <= P_14_1[28];
            mult_part_out01[291] <= P_8_5[35];
            mult_part_out01[292] <= P_6_7[22];
            mult_part_out01[293] <= P_14_1[31];
            mult_part_out01[294] <= P_7_6[31];
            mult_part_out01[295] <= P_7_7[8];
            mult_part_out01[296] <= P_3_9[29];
            mult_part_out01[297] <= P_13_2[28];
            mult_part_out01[298] <= P_6_7[28];
            mult_part_out01[299] <= P_7_6[36];
            mult_part_out01[300] <= P_4_8[40];
            mult_part_out01[301] <= P_4_9[17];
            mult_part_out01[302] <= P_9_6[5];
            mult_part_out01[303] <= P_7_7[16];
            mult_part_out01[304] <= P_13_2[35];
            mult_part_out01[305] <= P_15_2[2];
            mult_part_out01[306] <= P_9_5[33];
            mult_part_out01[307] <= P_9_6[10];
            mult_part_out01[308] <= P_6_8[14];
            mult_part_out01[309] <= P_4_9[25];
            mult_part_out01[310] <= P_6_8[16];
            mult_part_out01[311] <= P_14_3[1];
            mult_part_out01[312] <= P_11_5[5];
            mult_part_out01[313] <= P_5_9[12];
            mult_part_out01[314] <= P_12_4[14];
            mult_part_out01[315] <= P_7_8[4];
            mult_part_out01[316] <= P_12_3[40];
            mult_part_out01[317] <= P_10_6[3];
            mult_part_out01[318] <= P_10_6[4];
            mult_part_out01[319] <= P_12_4[19];
            mult_part_out01[320] <= P_7_7[33];
            mult_part_out01[321] <= P_3_10[30];
            mult_part_out01[322] <= P_7_7[35];
            mult_part_out01[323] <= P_13_4[6];
            mult_part_out01[324] <= P_13_3[31];
            mult_part_out01[325] <= P_9_6[28];
            mult_part_out01[326] <= P_5_10[1];
            mult_part_out01[327] <= P_9_6[30];
            mult_part_out01[328] <= P_8_7[24];
            mult_part_out01[329] <= P_13_3[36];
            mult_part_out01[330] <= P_10_6[16];
            mult_part_out01[331] <= P_10_6[17];
            mult_part_out01[332] <= P_8_8[4];
            mult_part_out01[333] <= P_11_5[26];
            mult_part_out01[334] <= P_4_10[26];
            mult_part_out01[335] <= P_14_3[25];
            mult_part_out01[336] <= P_14_4[2];
            mult_part_out01[337] <= P_15_3[10];
            mult_part_out01[338] <= P_7_8[27];
            mult_part_out01[339] <= P_9_7[18];
            mult_part_out01[340] <= P_6_9[22];
            mult_part_out01[341] <= P_6_9[23];
            mult_part_out01[342] <= P_8_8[14];
            mult_part_out01[343] <= P_14_4[9];
            mult_part_out01[344] <= P_13_5[3];
            mult_part_out01[345] <= P_13_4[28];
            mult_part_out01[346] <= P_10_7[8];
            mult_part_out01[347] <= P_11_6[16];
            mult_part_out01[348] <= P_8_8[20];
            mult_part_out01[349] <= P_9_7[28];
            mult_part_out01[350] <= P_9_7[29];
            mult_part_out01[351] <= P_13_5[10];
            mult_part_out01[352] <= P_12_6[4];
            mult_part_out01[353] <= P_12_5[29];
            mult_part_out01[354] <= P_13_4[37];
            mult_part_out01[355] <= P_5_10[30];
            mult_part_out01[356] <= P_14_4[22];
            mult_part_out01[357] <= P_11_6[26];
            mult_part_out01[358] <= P_11_7[3];
            mult_part_out01[359] <= P_8_8[31];
            mult_part_out01[360] <= P_8_8[32];
            mult_part_out01[361] <= P_8_9[9];
            mult_part_out01[362] <= P_11_7[7];
            mult_part_out01[363] <= P_12_6[15];
            mult_part_out01[364] <= P_15_4[13];
            mult_part_out01[365] <= P_9_8[20];
            mult_part_out01[366] <= P_7_9[31];
            mult_part_out01[367] <= P_11_7[12];
            mult_part_out01[368] <= P_10_7[30];
            mult_part_out01[369] <= P_11_7[14];
            mult_part_out01[370] <= P_13_5[29];
            mult_part_out01[371] <= P_10_8[9];
            mult_part_out01[372] <= P_9_8[27];
            mult_part_out01[373] <= P_8_9[21];
            mult_part_out01[374] <= P_6_10[32];
            mult_part_out01[375] <= P_11_7[20];
            mult_part_out01[376] <= P_13_5[35];
            mult_part_out01[377] <= P_10_7[39];
            mult_part_out01[378] <= P_10_7[40];
            mult_part_out01[379] <= P_12_7[7];
            mult_part_out01[380] <= P_9_9[11];
            mult_part_out01[381] <= P_7_10[22];
            mult_part_out01[382] <= P_11_7[27];
            mult_part_out01[383] <= P_9_8[38];
            mult_part_out01[384] <= P_10_8[22];
            mult_part_out01[385] <= P_14_6[3];
            mult_part_out01[386] <= P_9_9[17];
            mult_part_out01[387] <= P_11_7[32];
            mult_part_out01[388] <= P_10_8[26];
            mult_part_out01[389] <= P_9_9[20];
            mult_part_out01[390] <= P_8_10[14];
            mult_part_out01[391] <= P_11_8[12];
            mult_part_out01[392] <= P_14_6[10];
            mult_part_out01[393] <= P_14_5[35];
            mult_part_out01[394] <= P_10_8[32];
            mult_part_out01[395] <= P_10_9[9];
            mult_part_out01[396] <= P_13_6[31];
            mult_part_out01[397] <= P_8_10[21];
            mult_part_out01[398] <= P_12_8[2];
            mult_part_out01[399] <= P_9_10[6];
            mult_part_out01[400] <= P_10_9[14];
            mult_part_out01[401] <= P_9_9[32];
            mult_part_out01[402] <= P_8_10[26];
            mult_part_out01[403] <= P_11_8[24];
            mult_part_out01[404] <= P_13_6[39];
            mult_part_out01[405] <= P_8_10[29];
            mult_part_out01[406] <= P_12_8[10];
            mult_part_out01[407] <= P_10_9[21];
            mult_part_out01[408] <= P_11_9[5];
            mult_part_out01[409] <= P_14_6[27];
            mult_part_out01[410] <= P_10_9[24];
            mult_part_out01[411] <= P_14_7[5];
            mult_part_out01[412] <= P_14_6[30];
            mult_part_out01[413] <= P_13_7[24];
            mult_part_out01[414] <= P_11_9[11];
            mult_part_out01[415] <= P_11_8[36];
            mult_part_out01[416] <= P_14_6[34];
            mult_part_out01[417] <= P_11_9[14];
            mult_part_out01[418] <= P_10_10[8];
            mult_part_out01[419] <= P_12_8[23];
            mult_part_out01[420] <= P_10_10[10];
            mult_part_out01[421] <= P_9_10[28];
            mult_part_out01[422] <= P_13_7[33];
            mult_part_out01[423] <= P_10_9[37];
            mult_part_out01[424] <= P_10_10[14];
            mult_part_out01[425] <= P_9_10[32];
            mult_part_out01[426] <= P_13_7[37];
            mult_part_out01[427] <= P_14_7[21];
            mult_part_out01[428] <= P_13_7[39];
            mult_part_out01[429] <= P_12_9[9];
            mult_part_out01[430] <= P_14_8[0];
            mult_part_out01[431] <= P_15_7[8];
            mult_part_out01[432] <= P_11_9[29];
            mult_part_out01[433] <= P_11_10[6];
            mult_part_out01[434] <= P_13_8[21];
            mult_part_out01[435] <= P_13_8[22];
            mult_part_out01[436] <= P_12_8[40];
            mult_part_out01[437] <= P_15_7[14];
            mult_part_out01[438] <= P_13_8[25];
            mult_part_out01[439] <= P_13_8[26];
            mult_part_out01[440] <= P_14_8[10];
            mult_part_out01[441] <= P_11_9[38];
            mult_part_out01[442] <= P_13_9[5];
            mult_part_out01[443] <= P_15_7[20];
            mult_part_out01[444] <= P_12_10[0];
            mult_part_out01[445] <= P_15_7[22];
            mult_part_out01[446] <= P_13_9[9];
            mult_part_out01[447] <= P_15_8[0];
            mult_part_out01[448] <= P_13_8[35];
            mult_part_out01[449] <= P_13_9[12];
            mult_part_out01[450] <= P_13_9[13];
            mult_part_out01[451] <= P_13_9[14];
            mult_part_out01[452] <= P_13_9[15];
            mult_part_out01[453] <= P_15_8[6];
            mult_part_out01[454] <= P_11_10[27];
            mult_part_out01[455] <= P_11_10[28];
            mult_part_out01[456] <= P_14_8[26];
            mult_part_out01[457] <= P_13_9[20];
            mult_part_out01[458] <= P_14_9[4];
            mult_part_out01[459] <= P_15_8[12];
            mult_part_out01[460] <= P_15_8[13];
            mult_part_out01[461] <= P_13_10[0];
            mult_part_out01[462] <= P_14_9[8];
            mult_part_out01[463] <= P_12_10[19];
            mult_part_out01[464] <= P_14_9[10];
            mult_part_out01[465] <= P_15_8[18];
            mult_part_out01[466] <= P_14_8[36];
            mult_part_out01[467] <= P_14_9[13];
            mult_part_out01[468] <= P_12_10[24];
            mult_part_out01[469] <= P_13_9[32];
            mult_part_out01[470] <= P_14_9[16];
            mult_part_out01[471] <= P_13_10[10];
            mult_part_out01[472] <= P_15_9[1];
            mult_part_out01[473] <= P_13_10[12];
            mult_part_out01[474] <= P_15_9[3];
            mult_part_out01[475] <= P_13_10[14];
            mult_part_out01[476] <= P_12_10[32];
            mult_part_out01[477] <= P_14_9[23];
            mult_part_out01[478] <= P_13_10[17];
            mult_part_out01[479] <= P_15_9[8];
            mult_part_out01[480] <= P_14_10[2];
            mult_part_out01[481] <= P_14_10[3];
            mult_part_out01[482] <= P_13_10[21];
            mult_part_out01[483] <= P_13_10[22];
            mult_part_out01[484] <= P_14_9[30];
            mult_part_out01[485] <= P_13_10[24];
            mult_part_out01[486] <= P_14_10[8];
            mult_part_out01[487] <= P_14_10[9];
            mult_part_out01[488] <= P_14_10[10];
            mult_part_out01[489] <= P_15_9[18];
            mult_part_out01[490] <= P_14_9[36];
            mult_part_out01[491] <= P_15_9[20];
            mult_part_out01[492] <= P_14_9[38];
            mult_part_out01[493] <= P_13_10[32];
            mult_part_out01[494] <= P_14_10[16];
            mult_part_out01[495] <= P_14_10[17];
            mult_part_out01[496] <= P_14_10[18];
            mult_part_out01[497] <= P_15_10[2];
            mult_part_out01[498] <= P_14_10[20];
            mult_part_out01[499] <= P_15_10[4];
            mult_part_out01[500] <= P_14_10[22];
            mult_part_out01[501] <= P_15_10[6];
            mult_part_out01[502] <= P_14_10[24];
            mult_part_out01[503] <= P_15_10[8];
            mult_part_out01[504] <= P_15_10[9];
            mult_part_out01[505] <= P_15_10[10];
            mult_part_out01[506] <= P_14_10[28];
            mult_part_out01[507] <= P_15_10[12];
            mult_part_out01[508] <= P_14_10[30];
            mult_part_out01[509] <= P_15_10[14];
            mult_part_out01[510] <= P_15_10[15];

            mult_part_out02[24] <= P_0_1[0];
            mult_part_out02[25] <= P_1_0[8];
            mult_part_out02[26] <= P_1_0[9];
            mult_part_out02[27] <= P_0_0[27];
            mult_part_out02[28] <= P_1_0[11];
            mult_part_out02[29] <= P_1_0[12];
            mult_part_out02[30] <= P_0_0[30];
            mult_part_out02[31] <= P_0_1[7];
            mult_part_out02[32] <= P_1_0[15];
            mult_part_out02[33] <= P_0_1[9];
            mult_part_out02[34] <= P_1_0[17];
            mult_part_out02[35] <= P_1_0[18];
            mult_part_out02[36] <= P_0_0[36];
            mult_part_out02[37] <= P_0_1[13];
            mult_part_out02[38] <= P_1_0[21];
            mult_part_out02[39] <= P_0_0[39];
            mult_part_out02[40] <= P_0_0[40];
            mult_part_out02[41] <= P_1_0[24];
            mult_part_out02[42] <= P_0_1[18];
            mult_part_out02[43] <= P_1_0[26];
            mult_part_out02[44] <= P_1_0[27];
            mult_part_out02[45] <= P_1_1[4];
            mult_part_out02[46] <= P_1_0[29];
            mult_part_out02[47] <= P_2_0[13];
            mult_part_out02[48] <= P_0_1[24];
            mult_part_out02[49] <= P_1_1[8];
            mult_part_out02[50] <= P_0_2[2];
            mult_part_out02[51] <= P_0_1[27];
            mult_part_out02[52] <= P_2_0[18];
            mult_part_out02[53] <= P_1_1[12];
            mult_part_out02[54] <= P_2_0[20];
            mult_part_out02[55] <= P_0_1[31];
            mult_part_out02[56] <= P_3_0[5];
            mult_part_out02[57] <= P_0_2[9];
            mult_part_out02[58] <= P_1_1[17];
            mult_part_out02[59] <= P_3_0[8];
            mult_part_out02[60] <= P_0_1[36];
            mult_part_out02[61] <= P_0_2[13];
            mult_part_out02[62] <= P_1_1[21];
            mult_part_out02[63] <= P_2_0[29];
            mult_part_out02[64] <= P_2_1[6];
            mult_part_out02[65] <= P_2_0[31];
            mult_part_out02[66] <= P_1_2[1];
            mult_part_out02[67] <= P_2_1[9];
            mult_part_out02[68] <= P_4_0[0];
            mult_part_out02[69] <= P_3_0[18];
            mult_part_out02[70] <= P_2_0[36];
            mult_part_out02[71] <= P_4_0[3];
            mult_part_out02[72] <= P_2_1[14];
            mult_part_out02[73] <= P_0_3[1];
            mult_part_out02[74] <= P_3_0[23];
            mult_part_out02[75] <= P_4_0[7];
            mult_part_out02[76] <= P_2_1[18];
            mult_part_out02[77] <= P_1_1[36];
            mult_part_out02[78] <= P_1_1[37];
            mult_part_out02[79] <= P_4_0[11];
            mult_part_out02[80] <= P_3_1[5];
            mult_part_out02[81] <= P_0_3[9];
            mult_part_out02[82] <= P_3_1[7];
            mult_part_out02[83] <= P_2_1[25];
            mult_part_out02[84] <= P_3_1[9];
            mult_part_out02[85] <= P_2_2[3];
            mult_part_out02[86] <= P_3_1[11];
            mult_part_out02[87] <= P_4_0[19];
            mult_part_out02[88] <= P_4_0[20];
            mult_part_out02[89] <= P_0_3[17];
            mult_part_out02[90] <= P_3_1[15];
            mult_part_out02[91] <= P_5_0[6];
            mult_part_out02[92] <= P_2_1[34];
            mult_part_out02[93] <= P_4_1[1];
            mult_part_out02[94] <= P_1_2[29];
            mult_part_out02[95] <= P_0_3[23];
            mult_part_out02[96] <= P_0_4[0];
            mult_part_out02[97] <= P_1_2[32];
            mult_part_out02[98] <= P_4_0[30];
            mult_part_out02[99] <= P_5_0[14];
            mult_part_out02[100] <= P_0_4[4];
            mult_part_out02[101] <= P_2_2[19];
            mult_part_out02[102] <= P_1_3[13];
            mult_part_out02[103] <= P_0_3[31];
            mult_part_out02[104] <= P_4_0[36];
            mult_part_out02[105] <= P_5_0[20];
            mult_part_out02[106] <= P_4_0[38];
            mult_part_out02[107] <= P_4_1[15];
            mult_part_out02[108] <= P_0_3[36];
            mult_part_out02[109] <= P_0_4[13];
            mult_part_out02[110] <= P_1_3[21];
            mult_part_out02[111] <= P_4_1[19];
            mult_part_out02[112] <= P_0_3[40];
            mult_part_out02[113] <= P_6_0[11];
            mult_part_out02[114] <= P_2_2[32];
            mult_part_out02[115] <= P_1_4[2];
            mult_part_out02[116] <= P_5_1[7];
            mult_part_out02[117] <= P_5_0[32];
            mult_part_out02[118] <= P_4_1[26];
            mult_part_out02[119] <= P_4_2[3];
            mult_part_out02[120] <= P_2_2[38];
            mult_part_out02[121] <= P_1_4[8];
            mult_part_out02[122] <= P_6_0[20];
            mult_part_out02[123] <= P_0_4[27];
            mult_part_out02[124] <= P_0_5[4];
            mult_part_out02[125] <= P_4_1[33];
            mult_part_out02[126] <= P_0_4[30];
            mult_part_out02[127] <= P_6_0[25];
            mult_part_out02[128] <= P_0_5[8];
            mult_part_out02[129] <= P_2_3[23];
            mult_part_out02[130] <= P_2_3[24];
            mult_part_out02[131] <= P_5_1[22];
            mult_part_out02[132] <= P_2_3[26];
            mult_part_out02[133] <= P_0_5[13];
            mult_part_out02[134] <= P_3_3[11];
            mult_part_out02[135] <= P_2_3[29];
            mult_part_out02[136] <= P_6_1[10];
            mult_part_out02[137] <= P_7_0[18];
            mult_part_out02[138] <= P_5_1[29];
            mult_part_out02[139] <= P_6_1[13];
            mult_part_out02[140] <= P_3_3[17];
            mult_part_out02[141] <= P_4_2[25];
            mult_part_out02[142] <= P_0_5[22];
            mult_part_out02[143] <= P_5_1[34];
            mult_part_out02[144] <= P_0_5[24];
            mult_part_out02[145] <= P_1_5[8];
            mult_part_out02[146] <= P_1_5[9];
            mult_part_out02[147] <= P_2_4[17];
            mult_part_out02[148] <= P_8_0[12];
            mult_part_out02[149] <= P_4_2[33];
            mult_part_out02[150] <= P_1_4[37];
            mult_part_out02[151] <= P_0_6[7];
            mult_part_out02[152] <= P_7_0[33];
            mult_part_out02[153] <= P_1_4[40];
            mult_part_out02[154] <= P_8_0[18];
            mult_part_out02[155] <= P_4_2[39];
            mult_part_out02[156] <= P_2_4[26];
            mult_part_out02[157] <= P_6_2[7];
            mult_part_out02[158] <= P_0_6[14];
            mult_part_out02[159] <= P_9_0[6];
            mult_part_out02[160] <= P_5_2[27];
            mult_part_out02[161] <= P_9_0[8];
            mult_part_out02[162] <= P_9_0[9];
            mult_part_out02[163] <= P_3_3[40];
            mult_part_out02[164] <= P_4_4[0];
            mult_part_out02[165] <= P_7_1[22];
            mult_part_out02[166] <= P_1_6[5];
            mult_part_out02[167] <= P_5_3[10];
            mult_part_out02[168] <= P_5_3[11];
            mult_part_out02[169] <= P_7_1[26];
            mult_part_out02[170] <= P_4_4[6];
            mult_part_out02[171] <= P_5_2[38];
            mult_part_out02[172] <= P_0_6[28];
            mult_part_out02[173] <= P_1_5[36];
            mult_part_out02[174] <= P_7_2[7];
            mult_part_out02[175] <= P_1_6[14];
            mult_part_out02[176] <= P_4_4[12];
            mult_part_out02[177] <= P_0_7[9];
            mult_part_out02[178] <= P_8_1[18];
            mult_part_out02[179] <= P_3_5[8];
            mult_part_out02[180] <= P_4_3[40];
            mult_part_out02[181] <= P_6_3[7];
            mult_part_out02[182] <= P_6_3[8];
            mult_part_out02[183] <= P_8_1[23];
            mult_part_out02[184] <= P_8_1[24];
            mult_part_out02[185] <= P_5_3[28];
            mult_part_out02[186] <= P_7_2[19];
            mult_part_out02[187] <= P_1_6[26];
            mult_part_out02[188] <= P_4_4[24];
            mult_part_out02[189] <= P_9_1[12];
            mult_part_out02[190] <= P_9_0[37];
            mult_part_out02[191] <= P_8_1[31];
            mult_part_out02[192] <= P_2_6[14];
            mult_part_out02[193] <= P_8_2[9];
            mult_part_out02[194] <= P_8_2[10];
            mult_part_out02[195] <= P_10_1[1];
            mult_part_out02[196] <= P_0_7[28];
            mult_part_out02[197] <= P_3_5[26];
            mult_part_out02[198] <= P_0_7[30];
            mult_part_out02[199] <= P_7_2[32];
            mult_part_out02[200] <= P_10_0[30];
            mult_part_out02[201] <= P_10_0[31];
            mult_part_out02[202] <= P_2_7[0];
            mult_part_out02[203] <= P_8_2[19];
            mult_part_out02[204] <= P_4_5[16];
            mult_part_out02[205] <= P_2_6[27];
            mult_part_out02[206] <= P_5_4[25];
            mult_part_out02[207] <= P_12_0[3];
            mult_part_out02[208] <= P_0_8[16];
            mult_part_out02[209] <= P_4_5[21];
            mult_part_out02[210] <= P_12_0[6];
            mult_part_out02[211] <= P_10_1[17];
            mult_part_out02[212] <= P_1_7[27];
            mult_part_out02[213] <= P_4_6[1];
            mult_part_out02[214] <= P_9_1[37];
            mult_part_out02[215] <= P_1_8[6];
            mult_part_out02[216] <= P_9_1[39];
            mult_part_out02[217] <= P_8_3[9];
            mult_part_out02[218] <= P_0_9[2];
            mult_part_out02[219] <= P_12_0[15];
            mult_part_out02[220] <= P_0_9[4];
            mult_part_out02[221] <= P_8_2[37];
            mult_part_out02[222] <= P_11_0[35];
            mult_part_out02[223] <= P_0_9[7];
            mult_part_out02[224] <= P_0_8[32];
            mult_part_out02[225] <= P_8_3[17];
            mult_part_out02[226] <= P_10_2[8];
            mult_part_out02[227] <= P_2_7[25];
            mult_part_out02[228] <= P_0_8[36];
            mult_part_out02[229] <= P_7_4[14];
            mult_part_out02[230] <= P_5_6[1];
            mult_part_out02[231] <= P_9_2[30];
            mult_part_out02[232] <= P_12_1[4];
            mult_part_out02[233] <= P_1_9[0];
            mult_part_out02[234] <= P_12_1[6];
            mult_part_out02[235] <= P_9_2[34];
            mult_part_out02[236] <= P_4_6[24];
            mult_part_out02[237] <= P_6_5[15];
            mult_part_out02[238] <= P_1_9[5];
            mult_part_out02[239] <= P_5_5[34];
            mult_part_out02[240] <= P_13_0[19];
            mult_part_out02[241] <= P_3_7[22];
            mult_part_out02[242] <= P_7_5[3];
            mult_part_out02[243] <= P_12_0[39];
            mult_part_out02[244] <= P_4_6[32];
            mult_part_out02[245] <= P_7_4[30];
            mult_part_out02[246] <= P_10_3[4];
            mult_part_out02[247] <= P_1_8[38];
            mult_part_out02[248] <= P_0_10[8];
            mult_part_out02[249] <= P_9_4[0];
            mult_part_out02[250] <= P_6_5[28];
            mult_part_out02[251] <= P_11_1[40];
            mult_part_out02[252] <= P_11_2[17];
            mult_part_out02[253] <= P_7_4[38];
            mult_part_out02[254] <= P_3_8[11];
            mult_part_out02[255] <= P_12_2[3];
            mult_part_out02[256] <= P_7_5[17];
            mult_part_out02[257] <= P_12_1[29];
            mult_part_out02[258] <= P_7_5[19];
            mult_part_out02[259] <= P_11_2[24];
            mult_part_out02[260] <= P_0_10[20];
            mult_part_out02[261] <= P_6_6[15];
            mult_part_out02[262] <= P_0_10[22];
            mult_part_out02[263] <= P_3_8[20];
            mult_part_out02[264] <= P_14_0[26];
            mult_part_out02[265] <= P_11_3[6];
            mult_part_out02[266] <= P_5_6[37];
            mult_part_out02[267] <= P_0_10[27];
            mult_part_out02[268] <= P_1_10[11];
            mult_part_out02[269] <= P_7_5[30];
            mult_part_out02[270] <= P_4_7[34];
            mult_part_out02[271] <= P_3_8[28];
            mult_part_out02[272] <= P_0_10[32];
            mult_part_out02[273] <= P_13_2[4];
            mult_part_out02[274] <= P_12_2[22];
            mult_part_out02[275] <= P_2_9[25];
            mult_part_out02[276] <= P_3_8[33];
            mult_part_out02[277] <= P_5_8[0];
            mult_part_out02[278] <= P_5_8[1];
            mult_part_out02[279] <= P_6_6[33];
            mult_part_out02[280] <= P_11_3[21];
            mult_part_out02[281] <= P_3_8[38];
            mult_part_out02[282] <= P_7_6[19];
            mult_part_out02[283] <= P_10_4[17];
            mult_part_out02[284] <= P_1_10[27];
            mult_part_out02[285] <= P_4_9[1];
            mult_part_out02[286] <= P_1_10[29];
            mult_part_out02[287] <= P_8_6[7];
            mult_part_out02[288] <= P_5_7[35];
            mult_part_out02[289] <= P_15_1[10];
            mult_part_out02[290] <= P_4_8[30];
            mult_part_out02[291] <= P_14_2[5];
            mult_part_out02[292] <= P_14_2[6];
            mult_part_out02[293] <= P_13_2[24];
            mult_part_out02[294] <= P_13_3[1];
            mult_part_out02[295] <= P_3_10[4];
            mult_part_out02[296] <= P_6_8[2];
            mult_part_out02[297] <= P_9_6[0];
            mult_part_out02[298] <= P_3_9[31];
            mult_part_out02[299] <= P_14_2[13];
            mult_part_out02[300] <= P_3_9[33];
            mult_part_out02[301] <= P_6_8[7];
            mult_part_out02[302] <= P_14_2[16];
            mult_part_out02[303] <= P_10_5[13];
            mult_part_out02[304] <= P_8_7[0];
            mult_part_out02[305] <= P_3_9[38];
            mult_part_out02[306] <= P_12_3[30];
            mult_part_out02[307] <= P_14_2[21];
            mult_part_out02[308] <= P_11_5[1];
            mult_part_out02[309] <= P_6_7[39];
            mult_part_out02[310] <= P_4_10[2];
            mult_part_out02[311] <= P_5_8[34];
            mult_part_out02[312] <= P_3_10[21];
            mult_part_out02[313] <= P_12_3[37];
            mult_part_out02[314] <= P_11_5[7];
            mult_part_out02[315] <= P_8_7[11];
            mult_part_out02[316] <= P_8_6[36];
            mult_part_out02[317] <= P_11_5[10];
            mult_part_out02[318] <= P_8_7[14];
            mult_part_out02[319] <= P_13_3[26];
            mult_part_out02[320] <= P_4_9[36];
            mult_part_out02[321] <= P_11_5[14];
            mult_part_out02[322] <= P_9_6[25];
            mult_part_out02[323] <= P_14_2[37];
            mult_part_out02[324] <= P_14_2[38];
            mult_part_out02[325] <= P_12_4[25];
            mult_part_out02[326] <= P_6_9[8];
            mult_part_out02[327] <= P_12_4[27];
            mult_part_out02[328] <= P_8_8[0];
            mult_part_out02[329] <= P_12_4[29];
            mult_part_out02[330] <= P_9_6[33];
            mult_part_out02[331] <= P_14_3[21];
            mult_part_out02[332] <= P_10_6[18];
            mult_part_out02[333] <= P_6_9[15];
            mult_part_out02[334] <= P_8_8[6];
            mult_part_out02[335] <= P_5_9[34];
            mult_part_out02[336] <= P_8_7[32];
            mult_part_out02[337] <= P_4_10[29];
            mult_part_out02[338] <= P_11_6[7];
            mult_part_out02[339] <= P_4_10[31];
            mult_part_out02[340] <= P_10_6[26];
            mult_part_out02[341] <= P_5_10[16];
            mult_part_out02[342] <= P_6_10[0];
            mult_part_out02[343] <= P_15_3[16];
            mult_part_out02[344] <= P_10_7[6];
            mult_part_out02[345] <= P_14_3[35];
            mult_part_out02[346] <= P_11_5[39];
            mult_part_out02[347] <= P_12_5[23];
            mult_part_out02[348] <= P_10_7[10];
            mult_part_out02[349] <= P_5_10[24];
            mult_part_out02[350] <= P_13_4[33];
            mult_part_out02[351] <= P_9_7[30];
            mult_part_out02[352] <= P_13_5[11];
            mult_part_out02[353] <= P_6_9[35];
            mult_part_out02[354] <= P_15_4[3];
            mult_part_out02[355] <= P_13_5[14];
            mult_part_out02[356] <= P_10_7[18];
            mult_part_out02[357] <= P_11_7[2];
            mult_part_out02[358] <= P_9_8[13];
            mult_part_out02[359] <= P_13_5[18];
            mult_part_out02[360] <= P_9_7[39];
            mult_part_out02[361] <= P_9_8[16];
            mult_part_out02[362] <= P_10_7[24];
            mult_part_out02[363] <= P_8_8[35];
            mult_part_out02[364] <= P_9_8[19];
            mult_part_out02[365] <= P_7_9[30];
            mult_part_out02[366] <= P_8_8[38];
            mult_part_out02[367] <= P_14_4[33];
            mult_part_out02[368] <= P_14_4[34];
            mult_part_out02[369] <= P_10_8[7];
            mult_part_out02[370] <= P_10_8[8];
            mult_part_out02[371] <= P_10_7[33];
            mult_part_out02[372] <= P_13_5[31];
            mult_part_out02[373] <= P_7_9[38];
            mult_part_out02[374] <= P_8_9[22];
            mult_part_out02[375] <= P_14_5[17];
            mult_part_out02[376] <= P_8_9[24];
            mult_part_out02[377] <= P_11_7[22];
            mult_part_out02[378] <= P_10_8[16];
            mult_part_out02[379] <= P_8_10[3];
            mult_part_out02[380] <= P_11_7[25];
            mult_part_out02[381] <= P_13_5[40];
            mult_part_out02[382] <= P_9_9[13];
            mult_part_out02[383] <= P_10_8[21];
            mult_part_out02[384] <= P_13_6[19];
            mult_part_out02[385] <= P_11_8[6];
            mult_part_out02[386] <= P_12_7[14];
            mult_part_out02[387] <= P_8_9[35];
            mult_part_out02[388] <= P_12_7[16];
            mult_part_out02[389] <= P_14_5[31];
            mult_part_out02[390] <= P_13_7[1];
            mult_part_out02[391] <= P_8_10[15];
            mult_part_out02[392] <= P_13_6[27];
            mult_part_out02[393] <= P_10_8[31];
            mult_part_out02[394] <= P_15_5[19];
            mult_part_out02[395] <= P_9_10[2];
            mult_part_out02[396] <= P_12_7[24];
            mult_part_out02[397] <= P_13_7[8];
            mult_part_out02[398] <= P_13_6[33];
            mult_part_out02[399] <= P_10_8[37];
            mult_part_out02[400] <= P_13_6[35];
            mult_part_out02[401] <= P_11_8[22];
            mult_part_out02[402] <= P_11_8[23];
            mult_part_out02[403] <= P_12_8[7];
            mult_part_out02[404] <= P_14_6[22];
            mult_part_out02[405] <= P_9_9[36];
            mult_part_out02[406] <= P_14_6[24];
            mult_part_out02[407] <= P_14_7[1];
            mult_part_out02[408] <= P_8_10[32];
            mult_part_out02[409] <= P_15_6[10];
            mult_part_out02[410] <= P_13_7[21];
            mult_part_out02[411] <= P_11_9[8];
            mult_part_out02[412] <= P_10_10[2];
            mult_part_out02[413] <= P_11_8[34];
            mult_part_out02[414] <= P_11_8[35];
            mult_part_out02[415] <= P_13_7[26];
            mult_part_out02[416] <= P_13_7[27];
            mult_part_out02[417] <= P_13_7[28];
            mult_part_out02[418] <= P_14_7[12];
            mult_part_out02[419] <= P_15_6[20];
            mult_part_out02[420] <= P_12_9[0];
            mult_part_out02[421] <= P_12_9[1];
            mult_part_out02[422] <= P_12_9[2];
            mult_part_out02[423] <= P_13_7[34];
            mult_part_out02[424] <= P_12_8[28];
            mult_part_out02[425] <= P_13_8[12];
            mult_part_out02[426] <= P_13_8[13];
            mult_part_out02[427] <= P_13_8[14];
            mult_part_out02[428] <= P_12_9[8];
            mult_part_out02[429] <= P_14_7[23];
            mult_part_out02[430] <= P_11_9[27];
            mult_part_out02[431] <= P_14_8[1];
            mult_part_out02[432] <= P_10_10[22];
            mult_part_out02[433] <= P_15_7[10];
            mult_part_out02[434] <= P_14_7[28];
            mult_part_out02[435] <= P_11_9[32];
            mult_part_out02[436] <= P_11_10[9];
            mult_part_out02[437] <= P_13_9[0];
            mult_part_out02[438] <= P_11_9[35];
            mult_part_out02[439] <= P_11_9[36];
            mult_part_out02[440] <= P_13_8[27];
            mult_part_out02[441] <= P_12_9[21];
            mult_part_out02[442] <= P_15_7[19];
            mult_part_out02[443] <= P_13_8[30];
            mult_part_out02[444] <= P_15_7[21];
            mult_part_out02[445] <= P_11_10[18];
            mult_part_out02[446] <= P_11_10[19];
            mult_part_out02[447] <= P_15_7[24];
            mult_part_out02[448] <= P_12_10[4];
            mult_part_out02[449] <= P_12_9[29];
            mult_part_out02[450] <= P_11_10[23];
            mult_part_out02[451] <= P_12_9[31];
            mult_part_out02[452] <= P_14_8[22];
            mult_part_out02[453] <= P_12_10[9];
            mult_part_out02[454] <= P_12_10[10];
            mult_part_out02[455] <= P_12_9[35];
            mult_part_out02[456] <= P_12_10[12];
            mult_part_out02[457] <= P_11_10[30];
            mult_part_out02[458] <= P_15_8[11];
            mult_part_out02[459] <= P_11_10[32];
            mult_part_out02[460] <= P_13_9[23];
            mult_part_out02[461] <= P_14_9[7];
            mult_part_out02[462] <= P_15_8[15];
            mult_part_out02[463] <= P_13_9[26];
            mult_part_out02[464] <= P_12_10[20];
            mult_part_out02[465] <= P_13_9[28];
            mult_part_out02[466] <= P_13_9[29];
            mult_part_out02[467] <= P_13_9[30];
            mult_part_out02[468] <= P_13_9[31];
            mult_part_out02[469] <= P_15_8[22];
            mult_part_out02[470] <= P_13_9[33];
            mult_part_out02[471] <= P_15_9[0];
            mult_part_out02[472] <= P_13_10[11];
            mult_part_out02[473] <= P_14_9[19];
            mult_part_out02[474] <= P_13_9[37];
            mult_part_out02[475] <= P_15_9[4];
            mult_part_out02[476] <= P_13_9[39];
            mult_part_out02[477] <= P_13_10[16];
            mult_part_out02[478] <= P_14_9[24];
            mult_part_out02[479] <= P_14_9[25];
            mult_part_out02[480] <= P_15_9[9];
            mult_part_out02[481] <= P_15_9[10];
            mult_part_out02[482] <= P_14_10[4];
            mult_part_out02[483] <= P_14_10[5];
            mult_part_out02[484] <= P_13_10[23];
            mult_part_out02[485] <= P_14_9[31];
            mult_part_out02[486] <= P_14_9[32];
            mult_part_out02[487] <= P_15_9[16];
            mult_part_out02[488] <= P_13_10[27];
            mult_part_out02[489] <= P_13_10[28];
            mult_part_out02[490] <= P_15_9[19];
            mult_part_out02[491] <= P_13_10[30];
            mult_part_out02[492] <= P_13_10[31];
            mult_part_out02[493] <= P_15_9[22];
            mult_part_out02[494] <= P_14_9[40];
            mult_part_out02[495] <= P_15_9[24];

            mult_part_out03[34] <= P_0_1[10];
            mult_part_out03[35] <= P_0_1[11];
            mult_part_out03[36] <= P_0_1[12];
            mult_part_out03[37] <= P_0_0[37];
            mult_part_out03[38] <= P_2_0[4];
            mult_part_out03[39] <= P_0_1[15];
            mult_part_out03[40] <= P_2_0[6];
            mult_part_out03[41] <= P_2_0[7];
            mult_part_out03[42] <= P_2_0[8];
            mult_part_out03[43] <= P_2_0[9];
            mult_part_out03[44] <= P_1_1[3];
            mult_part_out03[45] <= P_2_0[11];
            mult_part_out03[46] <= P_1_1[5];
            mult_part_out03[47] <= P_1_1[6];
            mult_part_out03[48] <= P_1_0[31];
            mult_part_out03[49] <= P_0_1[25];
            mult_part_out03[50] <= P_1_0[33];
            mult_part_out03[51] <= P_0_2[3];
            mult_part_out03[52] <= P_3_0[1];
            mult_part_out03[53] <= P_1_0[36];
            mult_part_out03[54] <= P_3_0[3];
            mult_part_out03[55] <= P_1_0[38];
            mult_part_out03[56] <= P_0_1[32];
            mult_part_out03[57] <= P_1_1[16];
            mult_part_out03[58] <= P_2_1[0];
            mult_part_out03[59] <= P_2_1[1];
            mult_part_out03[60] <= P_1_1[19];
            mult_part_out03[61] <= P_2_0[27];
            mult_part_out03[62] <= P_3_0[11];
            mult_part_out03[63] <= P_3_0[12];
            mult_part_out03[64] <= P_2_0[30];
            mult_part_out03[65] <= P_1_2[0];
            mult_part_out03[66] <= P_2_0[32];
            mult_part_out03[67] <= P_1_1[26];
            mult_part_out03[68] <= P_3_0[17];
            mult_part_out03[69] <= P_1_1[28];
            mult_part_out03[70] <= P_1_2[5];
            mult_part_out03[71] <= P_2_1[13];
            mult_part_out03[72] <= P_3_0[21];
            mult_part_out03[73] <= P_0_2[25];
            mult_part_out03[74] <= P_1_2[9];
            mult_part_out03[75] <= P_1_2[10];
            mult_part_out03[76] <= P_0_3[4];
            mult_part_out03[77] <= P_0_2[29];
            mult_part_out03[78] <= P_1_2[13];
            mult_part_out03[79] <= P_0_3[7];
            mult_part_out03[80] <= P_0_2[32];
            mult_part_out03[81] <= P_1_1[40];
            mult_part_out03[82] <= P_2_1[24];
            mult_part_out03[83] <= P_0_3[11];
            mult_part_out03[84] <= P_2_1[26];
            mult_part_out03[85] <= P_1_2[20];
            mult_part_out03[86] <= P_0_2[38];
            mult_part_out03[87] <= P_3_1[12];
            mult_part_out03[88] <= P_3_1[13];
            mult_part_out03[89] <= P_3_1[14];
            mult_part_out03[90] <= P_0_3[18];
            mult_part_out03[91] <= P_4_0[23];
            mult_part_out03[92] <= P_3_1[17];
            mult_part_out03[93] <= P_5_0[8];
            mult_part_out03[94] <= P_3_1[19];
            mult_part_out03[95] <= P_4_1[3];
            mult_part_out03[96] <= P_4_1[4];
            mult_part_out03[97] <= P_5_0[12];
            mult_part_out03[98] <= P_2_2[16];
            mult_part_out03[99] <= P_3_2[0];
            mult_part_out03[100] <= P_1_3[11];
            mult_part_out03[101] <= P_0_3[29];
            mult_part_out03[102] <= P_2_2[20];
            mult_part_out03[103] <= P_1_2[38];
            mult_part_out03[104] <= P_3_1[29];
            mult_part_out03[105] <= P_4_0[37];
            mult_part_out03[106] <= P_6_0[4];
            mult_part_out03[107] <= P_1_3[18];
            mult_part_out03[108] <= P_1_3[19];
            mult_part_out03[109] <= P_5_1[0];
            mult_part_out03[110] <= P_5_0[25];
            mult_part_out03[111] <= P_2_2[29];
            mult_part_out03[112] <= P_5_0[27];
            mult_part_out03[113] <= P_5_1[4];
            mult_part_out03[114] <= P_6_0[12];
            mult_part_out03[115] <= P_2_2[33];
            mult_part_out03[116] <= P_5_0[31];
            mult_part_out03[117] <= P_1_3[28];
            mult_part_out03[118] <= P_5_1[9];
            mult_part_out03[119] <= P_2_2[37];
            mult_part_out03[120] <= P_1_4[7];
            mult_part_out03[121] <= P_2_2[39];
            mult_part_out03[122] <= P_0_4[26];
            mult_part_out03[123] <= P_3_2[24];
            mult_part_out03[124] <= P_7_0[5];
            mult_part_out03[125] <= P_7_0[6];
            mult_part_out03[126] <= P_7_0[7];
            mult_part_out03[127] <= P_0_5[7];
            mult_part_out03[128] <= P_2_3[22];
            mult_part_out03[129] <= P_4_1[37];
            mult_part_out03[130] <= P_3_2[31];
            mult_part_out03[131] <= P_1_4[18];
            mult_part_out03[132] <= P_4_2[16];
            mult_part_out03[133] <= P_3_3[10];
            mult_part_out03[134] <= P_6_1[8];
            mult_part_out03[135] <= P_1_4[22];
            mult_part_out03[136] <= P_5_1[27];
            mult_part_out03[137] <= P_3_2[38];
            mult_part_out03[138] <= P_2_4[8];
            mult_part_out03[139] <= P_5_1[30];
            mult_part_out03[140] <= P_0_5[20];
            mult_part_out03[141] <= P_1_4[28];
            mult_part_out03[142] <= P_3_3[19];
            mult_part_out03[143] <= P_3_3[20];
            mult_part_out03[144] <= P_2_4[14];
            mult_part_out03[145] <= P_4_3[5];
            mult_part_out03[146] <= P_7_0[27];
            mult_part_out03[147] <= P_3_4[0];
            mult_part_out03[148] <= P_3_4[1];
            mult_part_out03[149] <= P_4_3[9];
            mult_part_out03[150] <= P_4_2[34];
            mult_part_out03[151] <= P_2_4[21];
            mult_part_out03[152] <= P_1_5[15];
            mult_part_out03[153] <= P_5_2[20];
            mult_part_out03[154] <= P_6_1[28];
            mult_part_out03[155] <= P_6_1[29];
            mult_part_out03[156] <= P_8_0[20];
            mult_part_out03[157] <= P_3_4[10];
            mult_part_out03[158] <= P_6_2[8];
            mult_part_out03[159] <= P_6_2[9];
            mult_part_out03[160] <= P_3_3[37];
            mult_part_out03[161] <= P_1_5[24];
            mult_part_out03[162] <= P_8_0[26];
            mult_part_out03[163] <= P_8_0[27];
            mult_part_out03[164] <= P_8_0[28];
            mult_part_out03[165] <= P_5_2[32];
            mult_part_out03[166] <= P_8_0[30];
            mult_part_out03[167] <= P_0_6[23];
            mult_part_out03[168] <= P_3_4[21];
            mult_part_out03[169] <= P_7_2[2];
            mult_part_out03[170] <= P_5_2[37];
            mult_part_out03[171] <= P_1_5[34];
            mult_part_out03[172] <= P_3_4[25];
            mult_part_out03[173] <= P_4_4[9];
            mult_part_out03[174] <= P_4_3[34];
            mult_part_out03[175] <= P_9_0[22];
            mult_part_out03[176] <= P_7_1[33];
            mult_part_out03[177] <= P_8_1[17];
            mult_part_out03[178] <= P_4_4[14];
            mult_part_out03[179] <= P_0_6[35];
            mult_part_out03[180] <= P_3_5[9];
            mult_part_out03[181] <= P_7_1[38];
            mult_part_out03[182] <= P_3_5[11];
            mult_part_out03[183] <= P_6_2[33];
            mult_part_out03[184] <= P_3_5[13];
            mult_part_out03[185] <= P_6_2[35];
            mult_part_out03[186] <= P_6_3[12];
            mult_part_out03[187] <= P_5_3[30];
            mult_part_out03[188] <= P_5_4[7];
            mult_part_out03[189] <= P_8_1[29];
            mult_part_out03[190] <= P_10_0[20];
            mult_part_out03[191] <= P_2_6[13];
            mult_part_out03[192] <= P_8_2[8];
            mult_part_out03[193] <= P_7_2[26];
            mult_part_out03[194] <= P_6_3[20];
            mult_part_out03[195] <= P_6_3[21];
            mult_part_out03[196] <= P_10_1[2];
            mult_part_out03[197] <= P_9_1[20];
            mult_part_out03[198] <= P_7_2[31];
            mult_part_out03[199] <= P_1_6[38];
            mult_part_out03[200] <= P_1_6[39];
            mult_part_out03[201] <= P_6_4[3];
            mult_part_out03[202] <= P_6_4[4];
            mult_part_out03[203] <= P_7_3[12];
            mult_part_out03[204] <= P_6_4[6];
            mult_part_out03[205] <= P_3_5[34];
            mult_part_out03[206] <= P_3_6[11];
            mult_part_out03[207] <= P_10_1[13];
            mult_part_out03[208] <= P_6_4[10];
            mult_part_out03[209] <= P_12_0[5];
            mult_part_out03[210] <= P_9_1[33];
            mult_part_out03[211] <= P_9_2[10];
            mult_part_out03[212] <= P_5_4[31];
            mult_part_out03[213] <= P_12_0[9];
            mult_part_out03[214] <= P_6_4[16];
            mult_part_out03[215] <= P_11_1[4];
            mult_part_out03[216] <= P_0_9[0];
            mult_part_out03[217] <= P_4_6[5];
            mult_part_out03[218] <= P_10_2[0];
            mult_part_out03[219] <= P_11_0[32];
            mult_part_out03[220] <= P_2_7[18];
            mult_part_out03[221] <= P_13_0[0];
            mult_part_out03[222] <= P_7_3[31];
            mult_part_out03[223] <= P_6_4[25];
            mult_part_out03[224] <= P_10_1[30];
            mult_part_out03[225] <= P_0_8[33];
            mult_part_out03[226] <= P_4_6[14];
            mult_part_out03[227] <= P_8_3[19];
            mult_part_out03[228] <= P_3_6[33];
            mult_part_out03[229] <= P_6_5[7];
            mult_part_out03[230] <= P_13_0[9];
            mult_part_out03[231] <= P_3_7[12];
            mult_part_out03[232] <= P_3_6[37];
            mult_part_out03[233] <= P_6_4[35];
            mult_part_out03[234] <= P_1_9[1];
            mult_part_out03[235] <= P_8_3[27];
            mult_part_out03[236] <= P_13_0[15];
            mult_part_out03[237] <= P_0_9[21];
            mult_part_out03[238] <= P_5_6[9];
            mult_part_out03[239] <= P_8_4[7];
            mult_part_out03[240] <= P_5_5[35];
            mult_part_out03[241] <= P_12_1[13];
            mult_part_out03[242] <= P_12_0[38];
            mult_part_out03[243] <= P_11_2[8];
            mult_part_out03[244] <= P_10_2[26];
            mult_part_out03[245] <= P_9_3[20];
            mult_part_out03[246] <= P_14_0[8];
            mult_part_out03[247] <= P_2_8[21];
            mult_part_out03[248] <= P_3_7[29];
            mult_part_out03[249] <= P_11_1[38];
            mult_part_out03[250] <= P_11_2[15];
            mult_part_out03[251] <= P_8_4[19];
            mult_part_out03[252] <= P_7_5[13];
            mult_part_out03[253] <= P_2_9[3];
            mult_part_out03[254] <= P_10_3[12];
            mult_part_out03[255] <= P_14_0[17];
            mult_part_out03[256] <= P_5_6[27];
            mult_part_out03[257] <= P_2_8[31];
            mult_part_out03[258] <= P_14_0[20];
            mult_part_out03[259] <= P_1_9[26];
            mult_part_out03[260] <= P_6_6[14];
            mult_part_out03[261] <= P_12_1[33];
            mult_part_out03[262] <= P_5_7[9];
            mult_part_out03[263] <= P_11_3[4];
            mult_part_out03[264] <= P_7_5[25];
            mult_part_out03[265] <= P_15_0[10];
            mult_part_out03[266] <= P_3_8[23];
            mult_part_out03[267] <= P_9_4[18];
            mult_part_out03[268] <= P_12_1[40];
            mult_part_out03[269] <= P_11_3[10];
            mult_part_out03[270] <= P_2_9[20];
            mult_part_out03[271] <= P_1_9[38];
            mult_part_out03[272] <= P_9_4[23];
            mult_part_out03[273] <= P_3_8[30];
            mult_part_out03[274] <= P_14_0[36];
            mult_part_out03[275] <= P_1_10[18];
            mult_part_out03[276] <= P_12_2[24];
            mult_part_out03[277] <= P_9_5[4];
            mult_part_out03[278] <= P_9_4[29];
            mult_part_out03[279] <= P_9_5[6];
            mult_part_out03[280] <= P_6_7[10];
            mult_part_out03[281] <= P_1_10[24];
            mult_part_out03[282] <= P_13_1[37];
            mult_part_out03[283] <= P_12_3[7];
            mult_part_out03[284] <= P_15_1[5];
            mult_part_out03[285] <= P_10_4[19];
            mult_part_out03[286] <= P_7_6[23];
            mult_part_out03[287] <= P_10_4[21];
            mult_part_out03[288] <= P_2_9[38];
            mult_part_out03[289] <= P_9_4[40];
            mult_part_out03[290] <= P_10_5[0];
            mult_part_out03[291] <= P_5_8[14];
            mult_part_out03[292] <= P_2_10[18];
            mult_part_out03[293] <= P_2_10[19];
            mult_part_out03[294] <= P_10_4[28];
            mult_part_out03[295] <= P_10_5[5];
            mult_part_out03[296] <= P_11_4[13];
            mult_part_out03[297] <= P_9_5[24];
            mult_part_out03[298] <= P_11_3[39];
            mult_part_out03[299] <= P_3_9[32];
            mult_part_out03[300] <= P_9_5[27];
            mult_part_out03[301] <= P_3_9[34];
            mult_part_out03[302] <= P_12_3[26];
            mult_part_out03[303] <= P_12_3[27];
            mult_part_out03[304] <= P_5_9[3];
            mult_part_out03[305] <= P_10_5[15];
            mult_part_out03[306] <= P_12_4[6];
            mult_part_out03[307] <= P_11_4[24];
            mult_part_out03[308] <= P_12_4[8];
            mult_part_out03[309] <= P_11_4[26];
            mult_part_out03[310] <= P_11_5[3];
            mult_part_out03[311] <= P_4_9[27];
            mult_part_out03[312] <= P_5_8[35];
            mult_part_out03[313] <= P_4_10[5];
            mult_part_out03[314] <= P_3_10[23];
            mult_part_out03[315] <= P_4_10[7];
            mult_part_out03[316] <= P_10_6[2];
            mult_part_out03[317] <= P_7_7[30];
            mult_part_out03[318] <= P_4_9[34];
            mult_part_out03[319] <= P_13_4[2];
            mult_part_out03[320] <= P_10_5[30];
            mult_part_out03[321] <= P_5_9[20];
            mult_part_out03[322] <= P_4_9[38];
            mult_part_out03[323] <= P_12_4[23];
            mult_part_out03[324] <= P_5_9[23];
            mult_part_out03[325] <= P_6_9[7];
            mult_part_out03[326] <= P_10_5[36];
            mult_part_out03[327] <= P_8_7[23];
            mult_part_out03[328] <= P_15_3[1];
            mult_part_out03[329] <= P_9_7[8];
            mult_part_out03[330] <= P_15_3[3];
            mult_part_out03[331] <= P_12_5[7];
            mult_part_out03[332] <= P_5_9[31];
            mult_part_out03[333] <= P_13_4[16];
            mult_part_out03[334] <= P_6_8[40];
            mult_part_out03[335] <= P_5_10[10];
            mult_part_out03[336] <= P_5_9[35];
            mult_part_out03[337] <= P_7_9[2];
            mult_part_out03[338] <= P_9_7[17];
            mult_part_out03[339] <= P_6_9[21];
            mult_part_out03[340] <= P_5_10[15];
            mult_part_out03[341] <= P_12_5[17];
            mult_part_out03[342] <= P_5_10[17];
            mult_part_out03[343] <= P_5_10[18];
            mult_part_out03[344] <= P_14_4[10];
            mult_part_out03[345] <= P_6_9[27];
            mult_part_out03[346] <= P_14_4[12];
            mult_part_out03[347] <= P_13_4[30];
            mult_part_out03[348] <= P_5_10[23];
            mult_part_out03[349] <= P_8_8[21];
            mult_part_out03[350] <= P_12_6[2];
            mult_part_out03[351] <= P_15_3[24];
            mult_part_out03[352] <= P_8_9[0];
            mult_part_out03[353] <= P_13_4[36];
            mult_part_out03[354] <= P_11_6[23];
            mult_part_out03[355] <= P_13_4[38];
            mult_part_out03[356] <= P_8_8[28];
            mult_part_out03[357] <= P_7_9[22];
            mult_part_out03[358] <= P_6_9[40];
            mult_part_out03[359] <= P_9_7[38];
            mult_part_out03[360] <= P_14_5[2];
            mult_part_out03[361] <= P_11_6[30];
            mult_part_out03[362] <= P_8_8[34];
            mult_part_out03[363] <= P_10_8[1];
            mult_part_out03[364] <= P_12_6[16];
            mult_part_out03[365] <= P_10_8[3];
            mult_part_out03[366] <= P_13_5[25];
            mult_part_out03[367] <= P_9_8[22];
            mult_part_out03[368] <= P_15_4[17];
            mult_part_out03[369] <= P_12_6[21];
            mult_part_out03[370] <= P_9_9[1];
            mult_part_out03[371] <= P_14_4[37];
            mult_part_out03[372] <= P_8_9[20];
            mult_part_out03[373] <= P_12_6[25];
            mult_part_out03[374] <= P_13_6[9];
            mult_part_out03[375] <= P_8_9[23];
            mult_part_out03[376] <= P_12_7[4];
            mult_part_out03[377] <= P_12_6[29];
            mult_part_out03[378] <= P_9_8[33];
            mult_part_out03[379] <= P_13_5[38];
            mult_part_out03[380] <= P_15_5[5];
            mult_part_out03[381] <= P_9_8[36];
            mult_part_out03[382] <= P_15_5[7];
            mult_part_out03[383] <= P_11_8[4];
            mult_part_out03[384] <= P_7_10[25];
            mult_part_out03[385] <= P_12_6[37];
            mult_part_out03[386] <= P_11_7[31];
            mult_part_out03[387] <= P_12_6[39];
            mult_part_out03[388] <= P_14_5[30];
            mult_part_out03[389] <= P_10_9[3];
            mult_part_out03[390] <= P_8_9[38];
            mult_part_out03[391] <= P_12_7[19];
            mult_part_out03[392] <= P_8_10[16];
            mult_part_out03[393] <= P_11_8[14];
            mult_part_out03[394] <= P_12_7[22];
            mult_part_out03[395] <= P_14_5[37];
            mult_part_out03[396] <= P_10_8[34];
            mult_part_out03[397] <= P_13_6[32];
            mult_part_out03[398] <= P_11_8[19];
            mult_part_out03[399] <= P_10_9[13];
            mult_part_out03[400] <= P_14_6[18];
            mult_part_out03[401] <= P_9_10[8];
            mult_part_out03[402] <= P_14_6[20];
            mult_part_out03[403] <= P_14_6[21];
            mult_part_out03[404] <= P_8_10[28];
            mult_part_out03[405] <= P_9_10[12];
            mult_part_out03[406] <= P_9_10[13];
            mult_part_out03[407] <= P_8_10[31];
            mult_part_out03[408] <= P_13_7[19];
            mult_part_out03[409] <= P_12_7[37];
            mult_part_out03[410] <= P_12_8[14];
            mult_part_out03[411] <= P_14_6[29];
            mult_part_out03[412] <= P_15_6[13];
            mult_part_out03[413] <= P_10_10[3];
            mult_part_out03[414] <= P_10_10[4];
            mult_part_out03[415] <= P_14_6[33];
            mult_part_out03[416] <= P_14_7[10];
            mult_part_out03[417] <= P_12_8[21];
            mult_part_out03[418] <= P_13_7[29];
            mult_part_out03[419] <= P_10_10[9];
            mult_part_out03[420] <= P_11_9[17];
            mult_part_out03[421] <= P_11_9[18];
            mult_part_out03[422] <= P_10_10[12];
            mult_part_out03[423] <= P_9_10[30];
            mult_part_out03[424] <= P_15_7[1];
            mult_part_out03[425] <= P_11_9[22];
            mult_part_out03[426] <= P_10_10[16];
            mult_part_out03[427] <= P_13_7[38];
            mult_part_out03[428] <= P_11_9[25];
            mult_part_out03[429] <= P_11_9[26];
            mult_part_out03[430] <= P_11_10[3];
            mult_part_out03[431] <= P_11_10[4];
            mult_part_out03[432] <= P_12_8[36];
            mult_part_out03[433] <= P_14_7[27];
            mult_part_out03[434] <= P_11_9[31];
            mult_part_out03[435] <= P_10_10[25];
            mult_part_out03[436] <= P_13_8[23];
            mult_part_out03[437] <= P_14_7[31];
            mult_part_out03[438] <= P_11_10[11];
            mult_part_out03[439] <= P_15_7[16];
            mult_part_out03[440] <= P_13_9[3];
            mult_part_out03[441] <= P_14_8[11];
            mult_part_out03[442] <= P_11_9[39];
            mult_part_out03[443] <= P_14_8[13];
            mult_part_out03[444] <= P_13_8[31];
            mult_part_out03[445] <= P_12_9[25];
            mult_part_out03[446] <= P_14_8[16];
            mult_part_out03[447] <= P_13_9[10];
            mult_part_out03[448] <= P_11_10[21];
            mult_part_out03[449] <= P_14_8[19];
            mult_part_out03[450] <= P_12_10[6];
            mult_part_out03[451] <= P_13_8[38];
            mult_part_out03[452] <= P_13_8[39];
            mult_part_out03[453] <= P_13_9[16];
            mult_part_out03[454] <= P_14_8[24];
            mult_part_out03[455] <= P_14_9[1];
            mult_part_out03[456] <= P_12_9[36];
            mult_part_out03[457] <= P_14_9[3];
            mult_part_out03[458] <= P_12_10[14];
            mult_part_out03[459] <= P_14_9[5];
            mult_part_out03[460] <= P_14_9[6];
            mult_part_out03[461] <= P_15_8[14];
            mult_part_out03[462] <= P_13_9[25];
            mult_part_out03[463] <= P_15_8[16];
            mult_part_out03[464] <= P_14_8[34];
            mult_part_out03[465] <= P_14_9[11];
            mult_part_out03[466] <= P_14_9[12];
            mult_part_out03[467] <= P_12_10[23];
            mult_part_out03[468] <= P_14_8[38];
            mult_part_out03[469] <= P_12_10[25];
            mult_part_out03[470] <= P_14_8[40];
            mult_part_out03[471] <= P_15_8[24];
            mult_part_out03[472] <= P_13_9[35];
            mult_part_out03[473] <= P_13_9[36];
            mult_part_out03[474] <= P_12_10[30];
            mult_part_out03[475] <= P_14_9[21];
            mult_part_out03[476] <= P_15_9[5];
            mult_part_out03[477] <= P_15_9[6];
            mult_part_out03[478] <= P_15_9[7];
            mult_part_out03[479] <= P_13_10[18];
            mult_part_out03[480] <= P_13_10[19];
            mult_part_out03[481] <= P_13_10[20];
            mult_part_out03[482] <= P_14_9[28];
            mult_part_out03[483] <= P_15_9[12];
            mult_part_out03[484] <= P_15_9[13];
            mult_part_out03[485] <= P_14_10[7];
            mult_part_out03[486] <= P_15_9[15];
            mult_part_out03[487] <= P_14_9[33];
            mult_part_out03[488] <= P_14_9[34];
            mult_part_out03[489] <= P_14_9[35];
            mult_part_out03[490] <= P_13_10[29];
            mult_part_out03[491] <= P_14_10[13];
            mult_part_out03[492] <= P_15_9[21];
            mult_part_out03[493] <= P_14_9[39];

            mult_part_out04[48] <= P_2_0[14];
            mult_part_out04[49] <= P_2_0[15];
            mult_part_out04[50] <= P_0_1[26];
            mult_part_out04[51] <= P_2_0[17];
            mult_part_out04[52] <= P_0_1[28];
            mult_part_out04[53] <= P_0_2[5];
            mult_part_out04[54] <= P_0_1[30];
            mult_part_out04[55] <= P_0_2[7];
            mult_part_out04[56] <= P_1_1[15];
            mult_part_out04[57] <= P_0_1[33];
            mult_part_out04[58] <= P_0_1[34];
            mult_part_out04[59] <= P_1_1[18];
            mult_part_out04[60] <= P_3_0[9];
            mult_part_out04[61] <= P_0_1[37];
            mult_part_out04[62] <= P_2_1[4];
            mult_part_out04[63] <= P_2_1[5];
            mult_part_out04[64] <= P_0_2[16];
            mult_part_out04[65] <= P_1_1[24];
            mult_part_out04[66] <= P_0_2[18];
            mult_part_out04[67] <= P_1_2[2];
            mult_part_out04[68] <= P_2_1[10];
            mult_part_out04[69] <= P_4_0[1];
            mult_part_out04[70] <= P_3_0[19];
            mult_part_out04[71] <= P_1_2[6];
            mult_part_out04[72] <= P_4_0[4];
            mult_part_out04[73] <= P_2_1[15];
            mult_part_out04[74] <= P_4_0[6];
            mult_part_out04[75] <= P_2_1[17];
            mult_part_out04[76] <= P_3_0[25];
            mult_part_out04[77] <= P_3_0[26];
            mult_part_out04[78] <= P_3_0[27];
            mult_part_out04[79] <= P_1_2[14];
            mult_part_out04[80] <= P_1_2[15];
            mult_part_out04[81] <= P_4_0[13];
            mult_part_out04[82] <= P_0_3[10];
            mult_part_out04[83] <= P_4_0[15];
            mult_part_out04[84] <= P_1_2[19];
            mult_part_out04[85] <= P_4_0[17];
            mult_part_out04[86] <= P_2_2[4];
            mult_part_out04[87] <= P_2_1[29];
            mult_part_out04[88] <= P_0_3[16];
            mult_part_out04[89] <= P_2_1[31];
            mult_part_out04[90] <= P_1_2[25];
            mult_part_out04[91] <= P_1_2[26];
            mult_part_out04[92] <= P_1_2[27];
            mult_part_out04[93] <= P_0_3[21];
            mult_part_out04[94] <= P_1_3[5];
            mult_part_out04[95] <= P_1_2[30];
            mult_part_out04[96] <= P_5_0[11];
            mult_part_out04[97] <= P_0_4[1];
            mult_part_out04[98] <= P_0_3[26];
            mult_part_out04[99] <= P_1_2[34];
            mult_part_out04[100] <= P_5_0[15];
            mult_part_out04[101] <= P_3_2[2];
            mult_part_out04[102] <= P_0_4[6];
            mult_part_out04[103] <= P_4_1[11];
            mult_part_out04[104] <= P_6_0[2];
            mult_part_out04[105] <= P_6_0[3];
            mult_part_out04[106] <= P_3_1[31];
            mult_part_out04[107] <= P_3_1[32];
            mult_part_out04[108] <= P_5_0[23];
            mult_part_out04[109] <= P_2_2[27];
            mult_part_out04[110] <= P_6_0[8];
            mult_part_out04[111] <= P_6_0[9];
            mult_part_out04[112] <= P_6_0[10];
            mult_part_out04[113] <= P_4_1[21];
            mult_part_out04[114] <= P_3_1[39];
            mult_part_out04[115] <= P_6_0[13];
            mult_part_out04[116] <= P_6_0[14];
            mult_part_out04[117] <= P_2_2[35];
            mult_part_out04[118] <= P_5_0[33];
            mult_part_out04[119] <= P_0_4[23];
            mult_part_out04[120] <= P_0_4[24];
            mult_part_out04[121] <= P_4_1[29];
            mult_part_out04[122] <= P_4_1[30];
            mult_part_out04[123] <= P_1_4[10];
            mult_part_out04[124] <= P_1_4[11];
            mult_part_out04[125] <= P_5_0[40];
            mult_part_out04[126] <= P_1_4[13];
            mult_part_out04[127] <= P_7_0[8];
            mult_part_out04[128] <= P_3_2[29];
            mult_part_out04[129] <= P_7_0[10];
            mult_part_out04[130] <= P_6_0[28];
            mult_part_out04[131] <= P_3_2[32];
            mult_part_out04[132] <= P_7_0[13];
            mult_part_out04[133] <= P_5_1[24];
            mult_part_out04[134] <= P_0_4[38];
            mult_part_out04[135] <= P_0_5[15];
            mult_part_out04[136] <= P_7_0[17];
            mult_part_out04[137] <= P_3_3[14];
            mult_part_out04[138] <= P_6_1[12];
            mult_part_out04[139] <= P_6_0[37];
            mult_part_out04[140] <= P_1_4[27];
            mult_part_out04[141] <= P_5_1[32];
            mult_part_out04[142] <= P_8_0[6];
            mult_part_out04[143] <= P_7_0[24];
            mult_part_out04[144] <= P_7_0[25];
            mult_part_out04[145] <= P_0_5[25];
            mult_part_out04[146] <= P_4_2[30];
            mult_part_out04[147] <= P_1_5[10];
            mult_part_out04[148] <= P_5_2[15];
            mult_part_out04[149] <= P_2_4[19];
            mult_part_out04[150] <= P_5_2[17];
            mult_part_out04[151] <= P_3_4[4];
            mult_part_out04[152] <= P_3_4[5];
            mult_part_out04[153] <= P_4_2[37];
            mult_part_out04[154] <= P_3_4[7];
            mult_part_out04[155] <= P_3_4[8];
            mult_part_out04[156] <= P_3_4[9];
            mult_part_out04[157] <= P_0_6[13];
            mult_part_out04[158] <= P_3_4[11];
            mult_part_out04[159] <= P_1_5[22];
            mult_part_out04[160] <= P_1_5[23];
            mult_part_out04[161] <= P_4_3[21];
            mult_part_out04[162] <= P_4_3[22];
            mult_part_out04[163] <= P_5_3[6];
            mult_part_out04[164] <= P_6_2[14];
            mult_part_out04[165] <= P_9_0[12];
            mult_part_out04[166] <= P_5_2[33];
            mult_part_out04[167] <= P_1_5[30];
            mult_part_out04[168] <= P_0_7[0];
            mult_part_out04[169] <= P_5_2[36];
            mult_part_out04[170] <= P_3_4[23];
            mult_part_out04[171] <= P_4_3[31];
            mult_part_out04[172] <= P_1_5[35];
            mult_part_out04[173] <= P_5_2[40];
            mult_part_out04[174] <= P_3_4[27];
            mult_part_out04[175] <= P_1_5[38];
            mult_part_out04[176] <= P_6_3[2];
            mult_part_out04[177] <= P_4_4[13];
            mult_part_out04[178] <= P_7_1[35];
            mult_part_out04[179] <= P_1_6[18];
            mult_part_out04[180] <= P_7_1[37];
            mult_part_out04[181] <= P_9_1[4];
            mult_part_out04[182] <= P_1_6[21];
            mult_part_out04[183] <= P_3_4[36];
            mult_part_out04[184] <= P_5_4[3];
            mult_part_out04[185] <= P_1_7[0];
            mult_part_out04[186] <= P_2_5[32];
            mult_part_out04[187] <= P_2_5[33];
            mult_part_out04[188] <= P_8_2[4];
            mult_part_out04[189] <= P_4_5[1];
            mult_part_out04[190] <= P_7_2[23];
            mult_part_out04[191] <= P_4_5[3];
            mult_part_out04[192] <= P_2_5[38];
            mult_part_out04[193] <= P_1_7[8];
            mult_part_out04[194] <= P_1_7[9];
            mult_part_out04[195] <= P_9_1[18];
            mult_part_out04[196] <= P_5_4[15];
            mult_part_out04[197] <= P_0_8[5];
            mult_part_out04[198] <= P_10_0[28];
            mult_part_out04[199] <= P_10_0[29];
            mult_part_out04[200] <= P_3_5[29];
            mult_part_out04[201] <= P_10_1[7];
            mult_part_out04[202] <= P_10_0[32];
            mult_part_out04[203] <= P_3_6[8];
            mult_part_out04[204] <= P_0_7[36];
            mult_part_out04[205] <= P_7_3[14];
            mult_part_out04[206] <= P_8_2[22];
            mult_part_out04[207] <= P_7_2[40];
            mult_part_out04[208] <= P_8_3[0];
            mult_part_out04[209] <= P_8_3[1];
            mult_part_out04[210] <= P_10_1[16];
            mult_part_out04[211] <= P_1_8[2];
            mult_part_out04[212] <= P_9_1[35];
            mult_part_out04[213] <= P_5_4[32];
            mult_part_out04[214] <= P_1_8[5];
            mult_part_out04[215] <= P_12_0[11];
            mult_part_out04[216] <= P_0_8[24];
            mult_part_out04[217] <= P_11_1[6];
            mult_part_out04[218] <= P_1_8[9];
            mult_part_out04[219] <= P_7_3[28];
            mult_part_out04[220] <= P_1_7[35];
            mult_part_out04[221] <= P_1_8[12];
            mult_part_out04[222] <= P_12_0[18];
            mult_part_out04[223] <= P_7_4[8];
            mult_part_out04[224] <= P_2_7[22];
            mult_part_out04[225] <= P_5_5[20];
            mult_part_out04[226] <= P_5_5[21];
            mult_part_out04[227] <= P_0_8[35];
            mult_part_out04[228] <= P_9_2[27];
            mult_part_out04[229] <= P_10_2[11];
            mult_part_out04[230] <= P_8_3[22];
            mult_part_out04[231] <= P_6_4[33];
            mult_part_out04[232] <= P_8_3[24];
            mult_part_out04[233] <= P_10_2[15];
            mult_part_out04[234] <= P_9_3[9];
            mult_part_out04[235] <= P_11_1[24];
            mult_part_out04[236] <= P_10_2[18];
            mult_part_out04[237] <= P_1_8[28];
            mult_part_out04[238] <= P_2_7[36];
            mult_part_out04[239] <= P_4_6[27];
            mult_part_out04[240] <= P_10_2[22];
            mult_part_out04[241] <= P_9_2[40];
            mult_part_out04[242] <= P_14_0[4];
            mult_part_out04[243] <= P_14_0[5];
            mult_part_out04[244] <= P_1_9[11];
            mult_part_out04[245] <= P_13_1[0];
            mult_part_out04[246] <= P_1_9[13];
            mult_part_out04[247] <= P_8_3[39];
            mult_part_out04[248] <= P_11_2[13];
            mult_part_out04[249] <= P_2_8[23];
            mult_part_out04[250] <= P_8_4[18];
            mult_part_out04[251] <= P_9_4[2];
            mult_part_out04[252] <= P_10_3[10];
            mult_part_out04[253] <= P_13_0[32];
            mult_part_out04[254] <= P_11_2[19];
            mult_part_out04[255] <= P_15_0[0];
            mult_part_out04[256] <= P_12_2[4];
            mult_part_out04[257] <= P_6_5[35];
            mult_part_out04[258] <= P_10_2[40];
            mult_part_out04[259] <= P_15_0[4];
            mult_part_out04[260] <= P_5_7[7];
            mult_part_out04[261] <= P_10_3[19];
            mult_part_out04[262] <= P_14_0[24];
            mult_part_out04[263] <= P_5_7[10];
            mult_part_out04[264] <= P_5_7[11];
            mult_part_out04[265] <= P_0_10[25];
            mult_part_out04[266] <= P_7_5[27];
            mult_part_out04[267] <= P_12_1[39];
            mult_part_out04[268] <= P_13_1[23];
            mult_part_out04[269] <= P_8_4[37];
            mult_part_out04[270] <= P_13_1[25];
            mult_part_out04[271] <= P_2_9[21];
            mult_part_out04[272] <= P_8_4[40];
            mult_part_out04[273] <= P_9_4[24];
            mult_part_out04[274] <= P_9_5[1];
            mult_part_out04[275] <= P_3_8[32];
            mult_part_out04[276] <= P_7_5[37];
            mult_part_out04[277] <= P_11_3[18];
            mult_part_out04[278] <= P_12_2[26];
            mult_part_out04[279] <= P_3_8[36];
            mult_part_out04[280] <= P_5_7[27];
            mult_part_out04[281] <= P_4_8[21];
            mult_part_out04[282] <= P_9_4[33];
            mult_part_out04[283] <= P_7_6[20];
            mult_part_out04[284] <= P_11_4[1];
            mult_part_out04[285] <= P_11_4[2];
            mult_part_out04[286] <= P_6_7[16];
            mult_part_out04[287] <= P_12_3[11];
            mult_part_out04[288] <= P_4_8[28];
            mult_part_out04[289] <= P_5_8[12];
            mult_part_out04[290] <= P_7_7[3];
            mult_part_out04[291] <= P_12_3[15];
            mult_part_out04[292] <= P_11_3[33];
            mult_part_out04[293] <= P_8_5[37];
            mult_part_out04[294] <= P_4_8[34];
            mult_part_out04[295] <= P_15_1[16];
            mult_part_out04[296] <= P_14_2[10];
            mult_part_out04[297] <= P_7_6[34];
            mult_part_out04[298] <= P_10_5[8];
            mult_part_out04[299] <= P_9_6[2];
            mult_part_out04[300] <= P_3_10[9];
            mult_part_out04[301] <= P_9_5[28];
            mult_part_out04[302] <= P_13_2[33];
            mult_part_out04[303] <= P_2_10[29];
            mult_part_out04[304] <= P_12_3[28];
            mult_part_out04[305] <= P_9_6[8];
            mult_part_out04[306] <= P_10_5[16];
            mult_part_out04[307] <= P_5_9[6];
            mult_part_out04[308] <= P_7_7[21];
            mult_part_out04[309] <= P_15_2[6];
            mult_part_out04[310] <= P_11_4[27];
            mult_part_out04[311] <= P_6_8[17];
            mult_part_out04[312] <= P_14_3[2];
            mult_part_out04[313] <= P_11_4[30];
            mult_part_out04[314] <= P_13_3[21];
            mult_part_out04[315] <= P_11_5[8];
            mult_part_out04[316] <= P_4_10[8];
            mult_part_out04[317] <= P_8_6[37];
            mult_part_out04[318] <= P_4_10[10];
            mult_part_out04[319] <= P_11_5[12];
            mult_part_out04[320] <= P_6_8[26];
            mult_part_out04[321] <= P_8_7[17];
            mult_part_out04[322] <= P_9_7[1];
            mult_part_out04[323] <= P_10_5[33];
            mult_part_out04[324] <= P_15_2[21];
            mult_part_out04[325] <= P_5_10[0];
            mult_part_out04[326] <= P_7_8[15];
            mult_part_out04[327] <= P_7_7[40];
            mult_part_out04[328] <= P_6_8[34];
            mult_part_out04[329] <= P_12_5[5];
            mult_part_out04[330] <= P_9_7[9];
            mult_part_out04[331] <= P_5_10[6];
            mult_part_out04[332] <= P_13_3[39];
            mult_part_out04[333] <= P_7_8[22];
            mult_part_out04[334] <= P_13_4[17];
            mult_part_out04[335] <= P_9_6[38];
            mult_part_out04[336] <= P_15_3[9];
            mult_part_out04[337] <= P_6_9[19];
            mult_part_out04[338] <= P_7_9[3];
            mult_part_out04[339] <= P_8_8[11];
            mult_part_out04[340] <= P_14_4[6];
            mult_part_out04[341] <= P_14_4[7];
            mult_part_out04[342] <= P_11_6[11];
            mult_part_out04[343] <= P_12_5[19];
            mult_part_out04[344] <= P_11_6[13];
            mult_part_out04[345] <= P_8_8[17];
            mult_part_out04[346] <= P_15_3[19];
            mult_part_out04[347] <= P_5_10[22];
            mult_part_out04[348] <= P_12_6[0];
            mult_part_out04[349] <= P_9_8[4];
            mult_part_out04[350] <= P_14_4[16];
            mult_part_out04[351] <= P_8_8[23];
            mult_part_out04[352] <= P_7_9[17];
            mult_part_out04[353] <= P_14_4[19];
            mult_part_out04[354] <= P_7_9[19];
            mult_part_out04[355] <= P_12_5[31];
            mult_part_out04[356] <= P_6_10[14];
            mult_part_out04[357] <= P_13_5[16];
            mult_part_out04[358] <= P_8_8[30];
            mult_part_out04[359] <= P_6_10[17];
            mult_part_out04[360] <= P_14_4[26];
            mult_part_out04[361] <= P_6_10[19];
            mult_part_out04[362] <= P_7_10[3];
            mult_part_out04[363] <= P_13_5[22];
            mult_part_out04[364] <= P_7_10[5];
            mult_part_out04[365] <= P_11_6[34];
            mult_part_out04[366] <= P_14_4[32];
            mult_part_out04[367] <= P_8_9[15];
            mult_part_out04[368] <= P_11_6[37];
            mult_part_out04[369] <= P_13_6[4];
            mult_part_out04[370] <= P_14_5[12];
            mult_part_out04[371] <= P_11_7[16];
            mult_part_out04[372] <= P_14_4[38];
            mult_part_out04[373] <= P_13_6[8];
            mult_part_out04[374] <= P_12_7[2];
            mult_part_out04[375] <= P_12_6[27];
            mult_part_out04[376] <= P_7_10[17];
            mult_part_out04[377] <= P_13_6[12];
            mult_part_out04[378] <= P_8_9[26];
            mult_part_out04[379] <= P_11_7[24];
            mult_part_out04[380] <= P_14_5[22];
            mult_part_out04[381] <= P_9_9[12];
            mult_part_out04[382] <= P_10_8[20];
            mult_part_out04[383] <= P_15_5[8];
            mult_part_out04[384] <= P_12_7[12];
            mult_part_out04[385] <= P_14_5[27];
            mult_part_out04[386] <= P_10_9[0];
            mult_part_out04[387] <= P_14_5[29];
            mult_part_out04[388] <= P_15_5[13];
            mult_part_out04[389] <= P_11_7[34];
            mult_part_out04[390] <= P_12_7[18];
            mult_part_out04[391] <= P_7_10[32];
            mult_part_out04[392] <= P_14_5[34];
            mult_part_out04[393] <= P_9_10[0];
            mult_part_out04[394] <= P_11_8[15];
            mult_part_out04[395] <= P_12_7[23];
            mult_part_out04[396] <= P_8_10[20];
            mult_part_out04[397] <= P_10_9[11];
            mult_part_out04[398] <= P_10_9[12];
            mult_part_out04[399] <= P_15_6[0];
            mult_part_out04[400] <= P_13_7[11];
            mult_part_out04[401] <= P_10_9[15];
            mult_part_out04[402] <= P_10_8[40];
            mult_part_out04[403] <= P_12_7[31];
            mult_part_out04[404] <= P_11_8[25];
            mult_part_out04[405] <= P_13_7[16];
            mult_part_out04[406] <= P_11_9[3];
            mult_part_out04[407] <= P_9_9[38];
            mult_part_out04[408] <= P_12_8[12];
            mult_part_out04[409] <= P_9_9[40];
            mult_part_out04[410] <= P_12_7[38];
            mult_part_out04[411] <= P_9_10[18];
            mult_part_out04[412] <= P_9_10[19];
            mult_part_out04[413] <= P_14_7[7];
            mult_part_out04[414] <= P_13_7[25];
            mult_part_out04[415] <= P_15_6[16];
            mult_part_out04[416] <= P_10_9[30];
            mult_part_out04[417] <= P_14_6[35];
            mult_part_out04[418] <= P_13_8[5];
            mult_part_out04[419] <= P_14_6[37];
            mult_part_out04[420] <= P_9_10[27];
            mult_part_out04[421] <= P_13_8[8];
            mult_part_out04[422] <= P_14_6[40];
            mult_part_out04[423] <= P_12_9[3];
            mult_part_out04[424] <= P_11_9[21];
            mult_part_out04[425] <= P_10_9[39];
            mult_part_out04[426] <= P_12_9[6];
            mult_part_out04[427] <= P_11_10[0];
            mult_part_out04[428] <= P_13_8[15];
            mult_part_out04[429] <= P_13_8[16];
            mult_part_out04[430] <= P_13_8[17];
            mult_part_out04[431] <= P_13_8[18];
            mult_part_out04[432] <= P_14_8[2];
            mult_part_out04[433] <= P_13_8[20];
            mult_part_out04[434] <= P_15_7[11];
            mult_part_out04[435] <= P_14_8[5];
            mult_part_out04[436] <= P_12_9[16];
            mult_part_out04[437] <= P_11_9[34];
            mult_part_out04[438] <= P_12_9[18];
            mult_part_out04[439] <= P_14_7[33];
            mult_part_out04[440] <= P_15_7[17];
            mult_part_out04[441] <= P_15_7[18];
            mult_part_out04[442] <= P_11_10[15];
            mult_part_out04[443] <= P_12_9[23];
            mult_part_out04[444] <= P_14_7[38];
            mult_part_out04[445] <= P_14_8[15];
            mult_part_out04[446] <= P_13_8[33];
            mult_part_out04[447] <= P_12_9[27];
            mult_part_out04[448] <= P_13_9[11];
            mult_part_out04[449] <= P_13_8[36];
            mult_part_out04[450] <= P_12_9[30];
            mult_part_out04[451] <= P_15_8[4];
            mult_part_out04[452] <= P_12_9[32];
            mult_part_out04[453] <= P_12_9[33];
            mult_part_out04[454] <= P_13_9[17];
            mult_part_out04[455] <= P_12_10[11];
            mult_part_out04[456] <= P_11_10[29];
            mult_part_out04[457] <= P_12_9[37];
            mult_part_out04[458] <= P_11_10[31];
            mult_part_out04[459] <= P_13_9[22];
            mult_part_out04[460] <= P_14_8[30];
            mult_part_out04[461] <= P_12_10[17];
            mult_part_out04[462] <= P_13_10[1];
            mult_part_out04[463] <= P_14_8[33];
            mult_part_out04[464] <= P_13_9[27];
            mult_part_out04[465] <= P_12_10[21];
            mult_part_out04[466] <= P_12_10[22];
            mult_part_out04[467] <= P_13_10[6];
            mult_part_out04[468] <= P_15_8[21];
            mult_part_out04[469] <= P_14_9[15];
            mult_part_out04[470] <= P_15_8[23];
            mult_part_out04[471] <= P_13_9[34];
            mult_part_out04[472] <= P_12_10[28];
            mult_part_out04[473] <= P_15_9[2];
            mult_part_out04[474] <= P_14_9[20];
            mult_part_out04[475] <= P_13_9[38];
            mult_part_out04[476] <= P_14_9[22];

            mult_part_out05[51] <= P_3_0[0];
            mult_part_out05[52] <= P_1_1[11];
            mult_part_out05[53] <= P_2_0[19];
            mult_part_out05[54] <= P_1_1[13];
            mult_part_out05[55] <= P_2_0[21];
            mult_part_out05[56] <= P_1_0[39];
            mult_part_out05[57] <= P_1_0[40];
            mult_part_out05[58] <= P_2_0[24];
            mult_part_out05[59] <= P_0_1[35];
            mult_part_out05[60] <= P_2_1[2];
            mult_part_out05[61] <= P_3_0[10];
            mult_part_out05[62] <= P_0_2[14];
            mult_part_out05[63] <= P_1_1[22];
            mult_part_out05[64] <= P_1_1[23];
            mult_part_out05[65] <= P_0_2[17];
            mult_part_out05[66] <= P_2_1[8];
            mult_part_out05[67] <= P_0_2[19];
            mult_part_out05[68] <= P_0_2[20];
            mult_part_out05[69] <= P_1_2[4];
            mult_part_out05[70] <= P_1_1[29];
            mult_part_out05[71] <= P_3_0[20];
            mult_part_out05[72] <= P_1_2[7];
            mult_part_out05[73] <= P_1_1[32];
            mult_part_out05[74] <= P_2_0[40];
            mult_part_out05[75] <= P_0_3[3];
            mult_part_out05[76] <= P_1_2[11];
            mult_part_out05[77] <= P_4_0[9];
            mult_part_out05[78] <= P_3_1[3];
            mult_part_out05[79] <= P_2_1[21];
            mult_part_out05[80] <= P_1_1[39];
            mult_part_out05[81] <= P_3_1[6];
            mult_part_out05[82] <= P_0_2[34];
            mult_part_out05[83] <= P_0_2[35];
            mult_part_out05[84] <= P_3_0[33];
            mult_part_out05[85] <= P_0_3[13];
            mult_part_out05[86] <= P_1_2[21];
            mult_part_out05[87] <= P_0_3[15];
            mult_part_out05[88] <= P_2_1[30];
            mult_part_out05[89] <= P_1_3[0];
            mult_part_out05[90] <= P_5_0[5];
            mult_part_out05[91] <= P_3_1[16];
            mult_part_out05[92] <= P_1_3[3];
            mult_part_out05[93] <= P_4_0[25];
            mult_part_out05[94] <= P_2_2[12];
            mult_part_out05[95] <= P_2_2[13];
            mult_part_out05[96] <= P_3_1[21];
            mult_part_out05[97] <= P_3_1[22];
            mult_part_out05[98] <= P_5_0[13];
            mult_part_out05[99] <= P_3_1[24];
            mult_part_out05[100] <= P_2_2[18];
            mult_part_out05[101] <= P_1_3[12];
            mult_part_out05[102] <= P_6_0[0];
            mult_part_out05[103] <= P_3_1[28];
            mult_part_out05[104] <= P_5_0[19];
            mult_part_out05[105] <= P_2_2[23];
            mult_part_out05[106] <= P_1_3[17];
            mult_part_out05[107] <= P_4_0[39];
            mult_part_out05[108] <= P_4_1[16];
            mult_part_out05[109] <= P_1_3[20];
            mult_part_out05[110] <= P_4_1[18];
            mult_part_out05[111] <= P_0_4[15];
            mult_part_out05[112] <= P_1_3[23];
            mult_part_out05[113] <= P_5_0[28];
            mult_part_out05[114] <= P_5_0[29];
            mult_part_out05[115] <= P_2_3[9];
            mult_part_out05[116] <= P_3_2[17];
            mult_part_out05[117] <= P_0_4[21];
            mult_part_out05[118] <= P_4_2[2];
            mult_part_out05[119] <= P_1_4[6];
            mult_part_out05[120] <= P_7_0[1];
            mult_part_out05[121] <= P_2_3[15];
            mult_part_out05[122] <= P_1_4[9];
            mult_part_out05[123] <= P_5_1[14];
            mult_part_out05[124] <= P_2_3[18];
            mult_part_out05[125] <= P_2_3[19];
            mult_part_out05[126] <= P_2_3[20];
            mult_part_out05[127] <= P_0_4[31];
            mult_part_out05[128] <= P_7_0[9];
            mult_part_out05[129] <= P_3_2[30];
            mult_part_out05[130] <= P_6_1[4];
            mult_part_out05[131] <= P_0_5[11];
            mult_part_out05[132] <= P_0_4[36];
            mult_part_out05[133] <= P_3_2[34];
            mult_part_out05[134] <= P_4_2[18];
            mult_part_out05[135] <= P_5_1[26];
            mult_part_out05[136] <= P_0_5[16];
            mult_part_out05[137] <= P_8_0[1];
            mult_part_out05[138] <= P_7_0[19];
            mult_part_out05[139] <= P_1_5[2];
            mult_part_out05[140] <= P_4_3[0];
            mult_part_out05[141] <= P_1_5[4];
            mult_part_out05[142] <= P_2_3[36];
            mult_part_out05[143] <= P_7_1[0];
            mult_part_out05[144] <= P_0_6[0];
            mult_part_out05[145] <= P_2_4[15];
            mult_part_out05[146] <= P_2_4[16];
            mult_part_out05[147] <= P_3_3[24];
            mult_part_out05[148] <= P_7_0[29];
            mult_part_out05[149] <= P_0_6[5];
            mult_part_out05[150] <= P_3_3[27];
            mult_part_out05[151] <= P_4_3[11];
            mult_part_out05[152] <= P_7_1[9];
            mult_part_out05[153] <= P_2_4[23];
            mult_part_out05[154] <= P_7_1[11];
            mult_part_out05[155] <= P_8_0[19];
            mult_part_out05[156] <= P_0_6[12];
            mult_part_out05[157] <= P_5_3[0];
            mult_part_out05[158] <= P_2_4[28];
            mult_part_out05[159] <= P_4_3[19];
            mult_part_out05[160] <= P_8_0[24];
            mult_part_out05[161] <= P_8_0[25];
            mult_part_out05[162] <= P_2_5[8];
            mult_part_out05[163] <= P_8_1[3];
            mult_part_out05[164] <= P_1_5[27];
            mult_part_out05[165] <= P_5_3[8];
            mult_part_out05[166] <= P_7_1[23];
            mult_part_out05[167] <= P_4_3[27];
            mult_part_out05[168] <= P_2_4[38];
            mult_part_out05[169] <= P_0_7[1];
            mult_part_out05[170] <= P_9_0[17];
            mult_part_out05[171] <= P_3_4[24];
            mult_part_out05[172] <= P_2_5[18];
            mult_part_out05[173] <= P_4_3[33];
            mult_part_out05[174] <= P_4_4[10];
            mult_part_out05[175] <= P_2_5[21];
            mult_part_out05[176] <= P_0_6[32];
            mult_part_out05[177] <= P_6_3[3];
            mult_part_out05[178] <= P_1_6[17];
            mult_part_out05[179] <= P_0_7[11];
            mult_part_out05[180] <= P_0_6[36];
            mult_part_out05[181] <= P_2_5[27];
            mult_part_out05[182] <= P_5_3[25];
            mult_part_out05[183] <= P_1_6[22];
            mult_part_out05[184] <= P_6_3[10];
            mult_part_out05[185] <= P_1_6[24];
            mult_part_out05[186] <= P_1_7[1];
            mult_part_out05[187] <= P_1_7[2];
            mult_part_out05[188] <= P_0_7[20];
            mult_part_out05[189] <= P_2_6[11];
            mult_part_out05[190] <= P_0_7[22];
            mult_part_out05[191] <= P_4_4[27];
            mult_part_out05[192] <= P_9_0[39];
            mult_part_out05[193] <= P_2_5[39];
            mult_part_out05[194] <= P_3_5[23];
            mult_part_out05[195] <= P_2_6[17];
            mult_part_out05[196] <= P_8_2[12];
            mult_part_out05[197] <= P_1_6[36];
            mult_part_out05[198] <= P_8_2[14];
            mult_part_out05[199] <= P_3_5[28];
            mult_part_out05[200] <= P_6_3[26];
            mult_part_out05[201] <= P_7_3[10];
            mult_part_out05[202] <= P_7_3[11];
            mult_part_out05[203] <= P_6_3[29];
            mult_part_out05[204] <= P_4_4[40];
            mult_part_out05[205] <= P_6_4[7];
            mult_part_out05[206] <= P_10_0[36];
            mult_part_out05[207] <= P_3_6[12];
            mult_part_out05[208] <= P_11_0[21];
            mult_part_out05[209] <= P_2_6[31];
            mult_part_out05[210] <= P_7_3[19];
            mult_part_out05[211] <= P_1_7[26];
            mult_part_out05[212] <= P_6_3[38];
            mult_part_out05[213] <= P_8_2[29];
            mult_part_out05[214] <= P_0_8[22];
            mult_part_out05[215] <= P_5_5[10];
            mult_part_out05[216] <= P_5_4[35];
            mult_part_out05[217] <= P_10_1[23];
            mult_part_out05[218] <= P_0_8[26];
            mult_part_out05[219] <= P_8_3[11];
            mult_part_out05[220] <= P_6_4[22];
            mult_part_out05[221] <= P_8_3[13];
            mult_part_out05[222] <= P_1_7[37];
            mult_part_out05[223] <= P_4_6[11];
            mult_part_out05[224] <= P_1_8[15];
            mult_part_out05[225] <= P_10_1[31];
            mult_part_out05[226] <= P_0_8[34];
            mult_part_out05[227] <= P_6_4[29];
            mult_part_out05[228] <= P_8_3[20];
            mult_part_out05[229] <= P_9_3[4];
            mult_part_out05[230] <= P_11_1[19];
            mult_part_out05[231] <= P_4_6[19];
            mult_part_out05[232] <= P_0_9[16];
            mult_part_out05[233] <= P_6_5[11];
            mult_part_out05[234] <= P_1_8[25];
            mult_part_out05[235] <= P_3_7[16];
            mult_part_out05[236] <= P_12_1[8];
            mult_part_out05[237] <= P_4_7[1];
            mult_part_out05[238] <= P_6_4[40];
            mult_part_out05[239] <= P_7_5[0];
            mult_part_out05[240] <= P_7_5[1];
            mult_part_out05[241] <= P_10_2[23];
            mult_part_out05[242] <= P_1_8[33];
            mult_part_out05[243] <= P_10_2[25];
            mult_part_out05[244] <= P_12_0[40];
            mult_part_out05[245] <= P_5_5[40];
            mult_part_out05[246] <= P_4_6[34];
            mult_part_out05[247] <= P_11_1[36];
            mult_part_out05[248] <= P_6_6[2];
            mult_part_out05[249] <= P_3_8[6];
            mult_part_out05[250] <= P_9_4[1];
            mult_part_out05[251] <= P_0_9[35];
            mult_part_out05[252] <= P_9_4[3];
            mult_part_out05[253] <= P_14_0[15];
            mult_part_out05[254] <= P_6_5[32];
            mult_part_out05[255] <= P_7_4[40];
            mult_part_out05[256] <= P_9_3[31];
            mult_part_out05[257] <= P_8_4[25];
            mult_part_out05[258] <= P_4_7[22];
            mult_part_out05[259] <= P_8_4[27];
            mult_part_out05[260] <= P_10_3[18];
            mult_part_out05[261] <= P_11_2[26];
            mult_part_out05[262] <= P_9_3[37];
            mult_part_out05[263] <= P_7_5[24];
            mult_part_out05[264] <= P_12_2[12];
            mult_part_out05[265] <= P_11_2[30];
            mult_part_out05[266] <= P_4_8[6];
            mult_part_out05[267] <= P_1_9[34];
            mult_part_out05[268] <= P_14_0[30];
            mult_part_out05[269] <= P_10_3[27];
            mult_part_out05[270] <= P_10_4[4];
            mult_part_out05[271] <= P_10_4[5];
            mult_part_out05[272] <= P_7_6[9];
            mult_part_out05[273] <= P_15_0[18];
            mult_part_out05[274] <= P_10_4[8];
            mult_part_out05[275] <= P_9_4[26];
            mult_part_out05[276] <= P_2_9[26];
            mult_part_out05[277] <= P_13_1[32];
            mult_part_out05[278] <= P_4_8[18];
            mult_part_out05[279] <= P_4_8[19];
            mult_part_out05[280] <= P_8_5[24];
            mult_part_out05[281] <= P_5_8[4];
            mult_part_out05[282] <= P_6_6[36];
            mult_part_out05[283] <= P_13_1[38];
            mult_part_out05[284] <= P_9_5[11];
            mult_part_out05[285] <= P_5_8[8];
            mult_part_out05[286] <= P_11_4[3];
            mult_part_out05[287] <= P_12_2[35];
            mult_part_out05[288] <= P_10_4[22];
            mult_part_out05[289] <= P_2_10[15];
            mult_part_out05[290] <= P_15_1[11];
            mult_part_out05[291] <= P_6_7[21];
            mult_part_out05[292] <= P_8_6[12];
            mult_part_out05[293] <= P_6_7[23];
            mult_part_out05[294] <= P_6_7[24];
            mult_part_out05[295] <= P_10_4[29];
            mult_part_out05[296] <= P_3_10[5];
            mult_part_out05[297] <= P_2_10[23];
            mult_part_out05[298] <= P_13_3[5];
            mult_part_out05[299] <= P_4_9[15];
            mult_part_out05[300] <= P_6_8[6];
            mult_part_out05[301] <= P_3_10[10];
            mult_part_out05[302] <= P_3_9[35];
            mult_part_out05[303] <= P_15_2[0];
            mult_part_out05[304] <= P_4_9[20];
            mult_part_out05[305] <= P_10_4[39];
            mult_part_out05[306] <= P_4_9[22];
            mult_part_out05[307] <= P_15_2[4];
            mult_part_out05[308] <= P_15_2[5];
            mult_part_out05[309] <= P_12_3[33];
            mult_part_out05[310] <= P_14_2[24];
            mult_part_out05[311] <= P_12_3[35];
            mult_part_out05[312] <= P_9_5[39];
            mult_part_out05[313] <= P_6_8[19];
            mult_part_out05[314] <= P_6_8[20];
            mult_part_out05[315] <= P_12_4[15];
            mult_part_out05[316] <= P_10_5[26];
            mult_part_out05[317] <= P_12_4[17];
            mult_part_out05[318] <= P_13_4[1];
            mult_part_out05[319] <= P_9_6[22];
            mult_part_out05[320] <= P_3_10[29];
            mult_part_out05[321] <= P_6_9[3];
            mult_part_out05[322] <= P_3_10[31];
            mult_part_out05[323] <= P_7_8[12];
            mult_part_out05[324] <= P_6_8[30];
            mult_part_out05[325] <= P_5_9[24];
            mult_part_out05[326] <= P_5_9[25];
            mult_part_out05[327] <= P_9_7[6];
            mult_part_out05[328] <= P_13_4[11];
            mult_part_out05[329] <= P_4_10[21];
            mult_part_out05[330] <= P_6_9[12];
            mult_part_out05[331] <= P_13_3[38];
            mult_part_out05[332] <= P_5_10[7];
            mult_part_out05[333] <= P_4_10[25];
            mult_part_out05[334] <= P_10_6[20];
            mult_part_out05[335] <= P_12_4[35];
            mult_part_out05[336] <= P_7_8[25];
            mult_part_out05[337] <= P_12_5[13];
            mult_part_out05[338] <= P_5_10[13];
            mult_part_out05[339] <= P_5_10[14];
            mult_part_out05[340] <= P_10_7[2];
            mult_part_out05[341] <= P_8_7[37];
            mult_part_out05[342] <= P_11_5[35];
            mult_part_out05[343] <= P_10_6[29];
            mult_part_out05[344] <= P_15_3[17];
            mult_part_out05[345] <= P_12_5[21];
            mult_part_out05[346] <= P_9_7[25];
            mult_part_out05[347] <= P_13_5[6];
            mult_part_out05[348] <= P_14_4[14];
            mult_part_out05[349] <= P_7_9[14];
            mult_part_out05[350] <= P_14_3[40];
            mult_part_out05[351] <= P_9_8[6];
            mult_part_out05[352] <= P_9_8[7];
            mult_part_out05[353] <= P_6_10[11];
            mult_part_out05[354] <= P_5_10[29];
            mult_part_out05[355] <= P_15_4[4];
            mult_part_out05[356] <= P_12_5[32];
            mult_part_out05[357] <= P_10_7[19];
            mult_part_out05[358] <= P_10_7[20];
            mult_part_out05[359] <= P_11_7[4];
            mult_part_out05[360] <= P_11_7[5];
            mult_part_out05[361] <= P_13_5[20];
            mult_part_out05[362] <= P_14_5[4];
            mult_part_out05[363] <= P_8_9[11];
            mult_part_out05[364] <= P_12_5[40];
            mult_part_out05[365] <= P_12_6[17];
            mult_part_out05[366] <= P_6_10[24];
            mult_part_out05[367] <= P_13_6[2];
            mult_part_out05[368] <= P_7_9[33];
            mult_part_out05[369] <= P_7_9[34];
            mult_part_out05[370] <= P_15_4[19];
            mult_part_out05[371] <= P_15_4[20];
            mult_part_out05[372] <= P_12_7[0];
            mult_part_out05[373] <= P_9_8[28];
            mult_part_out05[374] <= P_12_6[26];
            mult_part_out05[375] <= P_13_6[10];
            mult_part_out05[376] <= P_10_8[14];
            mult_part_out05[377] <= P_13_5[36];
            mult_part_out05[378] <= P_8_10[2];
            mult_part_out05[379] <= P_8_9[27];
            mult_part_out05[380] <= P_10_8[18];
            mult_part_out05[381] <= P_10_8[19];
            mult_part_out05[382] <= P_9_8[37];
            mult_part_out05[383] <= P_14_5[25];
            mult_part_out05[384] <= P_11_7[29];
            mult_part_out05[385] <= P_7_10[26];
            mult_part_out05[386] <= P_10_8[24];
            mult_part_out05[387] <= P_8_10[11];
            mult_part_out05[388] <= P_13_6[23];
            mult_part_out05[389] <= P_12_7[17];
            mult_part_out05[390] <= P_13_6[25];
            mult_part_out05[391] <= P_10_8[29];
            mult_part_out05[392] <= P_15_5[17];
            mult_part_out05[393] <= P_13_6[28];
            mult_part_out05[394] <= P_11_7[39];
            mult_part_out05[395] <= P_11_8[16];
            mult_part_out05[396] <= P_9_10[3];
            mult_part_out05[397] <= P_14_5[39];
            mult_part_out05[398] <= P_13_7[9];
            mult_part_out05[399] <= P_15_5[24];
            mult_part_out05[400] <= P_8_10[24];
            mult_part_out05[401] <= P_13_6[36];
            mult_part_out05[402] <= P_10_9[16];
            mult_part_out05[403] <= P_15_6[4];
            mult_part_out05[404] <= P_9_9[35];
            mult_part_out05[405] <= P_13_6[40];
            mult_part_out05[406] <= P_14_7[0];
            mult_part_out05[407] <= P_9_10[14];
            mult_part_out05[408] <= P_9_9[39];
            mult_part_out05[409] <= P_13_7[20];
            mult_part_out05[410] <= P_10_10[0];
            mult_part_out05[411] <= P_11_8[32];
            mult_part_out05[412] <= P_11_8[33];
            mult_part_out05[413] <= P_11_9[10];
            mult_part_out05[414] <= P_15_6[15];
            mult_part_out05[415] <= P_10_10[5];
            mult_part_out05[416] <= P_10_10[6];
            mult_part_out05[417] <= P_9_10[24];
            mult_part_out05[418] <= P_10_9[32];
            mult_part_out05[419] <= P_9_10[26];
            mult_part_out05[420] <= P_12_8[24];
            mult_part_out05[421] <= P_12_8[25];
            mult_part_out05[422] <= P_13_8[9];
            mult_part_out05[423] <= P_10_10[13];
            mult_part_out05[424] <= P_9_10[31];
            mult_part_out05[425] <= P_14_7[19];
            mult_part_out05[426] <= P_15_7[3];
            mult_part_out05[427] <= P_15_7[4];
            mult_part_out05[428] <= P_14_7[22];
            mult_part_out05[429] <= P_12_8[33];
            mult_part_out05[430] <= P_14_7[24];
            mult_part_out05[431] <= P_12_8[35];
            mult_part_out05[432] <= P_15_7[9];
            mult_part_out05[433] <= P_12_9[13];
            mult_part_out05[434] <= P_14_8[4];
            mult_part_out05[435] <= P_12_8[39];
            mult_part_out05[436] <= P_10_10[26];
            mult_part_out05[437] <= P_12_9[17];
            mult_part_out05[438] <= P_15_7[15];
            mult_part_out05[439] <= P_12_9[19];
            mult_part_out05[440] <= P_14_7[34];
            mult_part_out05[441] <= P_14_7[35];
            mult_part_out05[442] <= P_14_8[12];
            mult_part_out05[443] <= P_14_7[37];
            mult_part_out05[444] <= P_12_9[24];
            mult_part_out05[445] <= P_13_8[32];
            mult_part_out05[446] <= P_14_7[40];
            mult_part_out05[447] <= P_11_10[20];
            mult_part_out05[448] <= P_12_9[28];
            mult_part_out05[449] <= P_11_10[22];
            mult_part_out05[450] <= P_14_8[20];
            mult_part_out05[451] <= P_12_10[7];
            mult_part_out05[452] <= P_15_8[5];
            mult_part_out05[453] <= P_14_8[23];
            mult_part_out05[454] <= P_12_9[34];
            mult_part_out05[455] <= P_13_9[18];
            mult_part_out05[456] <= P_15_8[9];
            mult_part_out05[457] <= P_14_8[27];
            mult_part_out05[458] <= P_14_8[28];
            mult_part_out05[459] <= P_14_8[29];
            mult_part_out05[460] <= P_12_9[40];
            mult_part_out05[461] <= P_13_9[24];
            mult_part_out05[462] <= P_14_8[32];
            mult_part_out05[463] <= P_13_10[2];
            mult_part_out05[464] <= P_13_10[3];
            mult_part_out05[465] <= P_13_10[4];
            mult_part_out05[466] <= P_13_10[5];
            mult_part_out05[467] <= P_14_8[37];
            mult_part_out05[468] <= P_14_9[14];
            mult_part_out05[469] <= P_13_10[8];
            mult_part_out05[470] <= P_12_10[26];
            mult_part_out05[471] <= P_14_9[17];

            mult_part_out06[68] <= P_2_0[34];
            mult_part_out06[69] <= P_2_0[35];
            mult_part_out06[70] <= P_0_2[22];
            mult_part_out06[71] <= P_2_0[37];
            mult_part_out06[72] <= P_0_2[24];
            mult_part_out06[73] <= P_4_0[5];
            mult_part_out06[74] <= P_2_1[16];
            mult_part_out06[75] <= P_0_2[27];
            mult_part_out06[76] <= P_3_1[1];
            mult_part_out06[77] <= P_3_1[2];
            mult_part_out06[78] <= P_4_0[10];
            mult_part_out06[79] <= P_3_0[28];
            mult_part_out06[80] <= P_4_0[12];
            mult_part_out06[81] <= P_2_1[23];
            mult_part_out06[82] <= P_1_2[17];
            mult_part_out06[83] <= P_1_2[18];
            mult_part_out06[84] <= P_2_2[2];
            mult_part_out06[85] <= P_3_1[10];
            mult_part_out06[86] <= P_3_0[35];
            mult_part_out06[87] <= P_0_2[39];
            mult_part_out06[88] <= P_5_0[3];
            mult_part_out06[89] <= P_1_2[24];
            mult_part_out06[90] <= P_2_1[32];
            mult_part_out06[91] <= P_2_1[33];
            mult_part_out06[92] <= P_0_3[20];
            mult_part_out06[93] <= P_1_3[4];
            mult_part_out06[94] <= P_4_0[26];
            mult_part_out06[95] <= P_2_1[37];
            mult_part_out06[96] <= P_1_3[7];
            mult_part_out06[97] <= P_2_2[15];
            mult_part_out06[98] <= P_3_1[23];
            mult_part_out06[99] <= P_1_3[10];
            mult_part_out06[100] <= P_3_2[1];
            mult_part_out06[101] <= P_4_0[33];
            mult_part_out06[102] <= P_5_0[17];
            mult_part_out06[103] <= P_1_3[14];
            mult_part_out06[104] <= P_1_3[15];
            mult_part_out06[105] <= P_3_2[6];
            mult_part_out06[106] <= P_2_2[24];
            mult_part_out06[107] <= P_2_2[25];
            mult_part_out06[108] <= P_2_3[2];
            mult_part_out06[109] <= P_5_0[24];
            mult_part_out06[110] <= P_3_1[35];
            mult_part_out06[111] <= P_3_2[12];
            mult_part_out06[112] <= P_3_1[37];
            mult_part_out06[113] <= P_1_3[24];
            mult_part_out06[114] <= P_4_1[22];
            mult_part_out06[115] <= P_1_3[26];
            mult_part_out06[116] <= P_0_4[20];
            mult_part_out06[117] <= P_1_4[4];
            mult_part_out06[118] <= P_1_4[5];
            mult_part_out06[119] <= P_6_0[17];
            mult_part_out06[120] <= P_4_1[28];
            mult_part_out06[121] <= P_4_2[5];
            mult_part_out06[122] <= P_5_0[37];
            mult_part_out06[123] <= P_6_0[21];
            mult_part_out06[124] <= P_4_2[8];
            mult_part_out06[125] <= P_0_5[5];
            mult_part_out06[126] <= P_4_2[10];
            mult_part_out06[127] <= P_3_2[28];
            mult_part_out06[128] <= P_1_3[39];
            mult_part_out06[129] <= P_0_4[33];
            mult_part_out06[130] <= P_2_4[0];
            mult_part_out06[131] <= P_6_0[29];
            mult_part_out06[132] <= P_1_4[19];
            mult_part_out06[133] <= P_6_1[7];
            mult_part_out06[134] <= P_2_4[4];
            mult_part_out06[135] <= P_5_2[2];
            mult_part_out06[136] <= P_3_2[37];
            mult_part_out06[137] <= P_6_1[11];
            mult_part_out06[138] <= P_5_2[5];
            mult_part_out06[139] <= P_5_2[6];
            mult_part_out06[140] <= P_8_0[4];
            mult_part_out06[141] <= P_6_0[39];
            mult_part_out06[142] <= P_2_4[12];
            mult_part_out06[143] <= P_1_5[6];
            mult_part_out06[144] <= P_8_0[8];
            mult_part_out06[145] <= P_8_0[9];
            mult_part_out06[146] <= P_0_5[26];
            mult_part_out06[147] <= P_4_2[31];
            mult_part_out06[148] <= P_6_1[22];
            mult_part_out06[149] <= P_3_4[2];
            mult_part_out06[150] <= P_6_1[24];
            mult_part_out06[151] <= P_4_2[35];
            mult_part_out06[152] <= P_5_2[19];
            mult_part_out06[153] <= P_3_4[6];
            mult_part_out06[154] <= P_2_5[0];
            mult_part_out06[155] <= P_9_0[2];
            mult_part_out06[156] <= P_7_0[37];
            mult_part_out06[157] <= P_2_5[3];
            mult_part_out06[158] <= P_7_0[39];
            mult_part_out06[159] <= P_8_0[23];
            mult_part_out06[160] <= P_0_5[40];
            mult_part_out06[161] <= P_3_4[14];
            mult_part_out06[162] <= P_5_3[5];
            mult_part_out06[163] <= P_2_5[9];
            mult_part_out06[164] <= P_5_2[31];
            mult_part_out06[165] <= P_4_3[25];
            mult_part_out06[166] <= P_1_5[29];
            mult_part_out06[167] <= P_2_4[37];
            mult_part_out06[168] <= P_4_3[28];
            mult_part_out06[169] <= P_8_1[9];
            mult_part_out06[170] <= P_0_7[2];
            mult_part_out06[171] <= P_0_7[3];
            mult_part_out06[172] <= P_10_0[2];
            mult_part_out06[173] <= P_8_0[37];
            mult_part_out06[174] <= P_3_5[3];
            mult_part_out06[175] <= P_5_3[18];
            mult_part_out06[176] <= P_3_4[29];
            mult_part_out06[177] <= P_3_4[30];
            mult_part_out06[178] <= P_0_7[10];
            mult_part_out06[179] <= P_2_5[25];
            mult_part_out06[180] <= P_7_2[13];
            mult_part_out06[181] <= P_6_2[31];
            mult_part_out06[182] <= P_3_4[35];
            mult_part_out06[183] <= P_7_1[40];
            mult_part_out06[184] <= P_0_6[40];
            mult_part_out06[185] <= P_3_4[38];
            mult_part_out06[186] <= P_3_5[15];
            mult_part_out06[187] <= P_10_0[17];
            mult_part_out06[188] <= P_10_0[18];
            mult_part_out06[189] <= P_5_4[8];
            mult_part_out06[190] <= P_4_4[26];
            mult_part_out06[191] <= P_7_2[24];
            mult_part_out06[192] <= P_10_0[22];
            mult_part_out06[193] <= P_9_1[16];
            mult_part_out06[194] <= P_2_6[16];
            mult_part_out06[195] <= P_7_2[28];
            mult_part_out06[196] <= P_8_1[36];
            mult_part_out06[197] <= P_10_0[27];
            mult_part_out06[198] <= P_8_1[38];
            mult_part_out06[199] <= P_1_7[14];
            mult_part_out06[200] <= P_6_4[2];
            mult_part_out06[201] <= P_9_1[24];
            mult_part_out06[202] <= P_1_7[17];
            mult_part_out06[203] <= P_6_4[5];
            mult_part_out06[204] <= P_5_4[23];
            mult_part_out06[205] <= P_4_5[17];
            mult_part_out06[206] <= P_9_2[5];
            mult_part_out06[207] <= P_5_4[26];
            mult_part_out06[208] <= P_2_7[6];
            mult_part_out06[209] <= P_7_3[18];
            mult_part_out06[210] <= P_10_0[40];
            mult_part_out06[211] <= P_5_5[6];
            mult_part_out06[212] <= P_5_5[7];
            mult_part_out06[213] <= P_8_3[5];
            mult_part_out06[214] <= P_9_2[13];
            mult_part_out06[215] <= P_10_1[21];
            mult_part_out06[216] <= P_8_3[8];
            mult_part_out06[217] <= P_0_9[1];
            mult_part_out06[218] <= P_7_4[3];
            mult_part_out06[219] <= P_9_2[18];
            mult_part_out06[220] <= P_4_6[8];
            mult_part_out06[221] <= P_7_3[30];
            mult_part_out06[222] <= P_4_5[34];
            mult_part_out06[223] <= P_8_2[39];
            mult_part_out06[224] <= P_13_0[3];
            mult_part_out06[225] <= P_2_7[23];
            mult_part_out06[226] <= P_10_1[32];
            mult_part_out06[227] <= P_0_9[11];
            mult_part_out06[228] <= P_11_1[17];
            mult_part_out06[229] <= P_10_1[35];
            mult_part_out06[230] <= P_6_5[8];
            mult_part_out06[231] <= P_0_8[39];
            mult_part_out06[232] <= P_7_4[17];
            mult_part_out06[233] <= P_7_4[18];
            mult_part_out06[234] <= P_8_3[26];
            mult_part_out06[235] <= P_6_5[13];
            mult_part_out06[236] <= P_11_2[1];
            mult_part_out06[237] <= P_2_8[11];
            mult_part_out06[238] <= P_11_2[3];
            mult_part_out06[239] <= P_1_9[6];
            mult_part_out06[240] <= P_2_8[14];
            mult_part_out06[241] <= P_2_8[15];
            mult_part_out06[242] <= P_8_3[34];
            mult_part_out06[243] <= P_1_8[34];
            mult_part_out06[244] <= P_8_4[12];
            mult_part_out06[245] <= P_12_1[17];
            mult_part_out06[246] <= P_4_7[10];
            mult_part_out06[247] <= P_3_8[4];
            mult_part_out06[248] <= P_8_4[16];
            mult_part_out06[249] <= P_4_7[13];
            mult_part_out06[250] <= P_5_6[21];
            mult_part_out06[251] <= P_13_1[6];
            mult_part_out06[252] <= P_13_0[31];
            mult_part_out06[253] <= P_0_10[13];
            mult_part_out06[254] <= P_5_7[1];
            mult_part_out06[255] <= P_3_7[36];
            mult_part_out06[256] <= P_4_7[20];
            mult_part_out06[257] <= P_0_10[17];
            mult_part_out06[258] <= P_1_9[25];
            mult_part_out06[259] <= P_10_3[17];
            mult_part_out06[260] <= P_8_5[4];
            mult_part_out06[261] <= P_5_7[8];
            mult_part_out06[262] <= P_12_1[34];
            mult_part_out06[263] <= P_2_8[37];
            mult_part_out06[264] <= P_10_3[22];
            mult_part_out06[265] <= P_13_1[20];
            mult_part_out06[266] <= P_5_7[13];
            mult_part_out06[267] <= P_2_9[17];
            mult_part_out06[268] <= P_5_6[39];
            mult_part_out06[269] <= P_0_10[29];
            mult_part_out06[270] <= P_3_8[27];
            mult_part_out06[271] <= P_11_2[36];
            mult_part_out06[272] <= P_1_9[39];
            mult_part_out06[273] <= P_6_6[27];
            mult_part_out06[274] <= P_6_7[4];
            mult_part_out06[275] <= P_7_5[36];
            mult_part_out06[276] <= P_10_4[10];
            mult_part_out06[277] <= P_6_6[31];
            mult_part_out06[278] <= P_9_5[5];
            mult_part_out06[279] <= P_11_3[20];
            mult_part_out06[280] <= P_8_6[0];
            mult_part_out06[281] <= P_14_1[19];
            mult_part_out06[282] <= P_8_5[26];
            mult_part_out06[283] <= P_5_7[30];
            mult_part_out06[284] <= P_12_2[32];
            mult_part_out06[285] <= P_1_10[28];
            mult_part_out06[286] <= P_11_3[27];
            mult_part_out06[287] <= P_11_4[4];
            mult_part_out06[288] <= P_7_7[1];
            mult_part_out06[289] <= P_12_3[13];
            mult_part_out06[290] <= P_8_5[34];
            mult_part_out06[291] <= P_4_8[31];
            mult_part_out06[292] <= P_7_6[29];
            mult_part_out06[293] <= P_9_5[20];
            mult_part_out06[294] <= P_2_10[20];
            mult_part_out06[295] <= P_8_5[39];
            mult_part_out06[296] <= P_12_3[20];
            mult_part_out06[297] <= P_14_1[35];
            mult_part_out06[298] <= P_3_10[7];
            mult_part_out06[299] <= P_10_4[33];
            mult_part_out06[300] <= P_10_4[34];
            mult_part_out06[301] <= P_14_1[39];
            mult_part_out06[302] <= P_8_6[22];
            mult_part_out06[303] <= P_7_6[40];
            mult_part_out06[304] <= P_6_8[10];
            mult_part_out06[305] <= P_7_7[18];
            mult_part_out06[306] <= P_15_2[3];
            mult_part_out06[307] <= P_13_2[38];
            mult_part_out06[308] <= P_4_10[0];
            mult_part_out06[309] <= P_12_4[9];
            mult_part_out06[310] <= P_7_7[23];
            mult_part_out06[311] <= P_7_8[0];
            mult_part_out06[312] <= P_4_9[28];
            mult_part_out06[313] <= P_7_8[2];
            mult_part_out06[314] <= P_5_8[37];
            mult_part_out06[315] <= P_10_5[25];
            mult_part_out06[316] <= P_13_3[23];
            mult_part_out06[317] <= P_9_6[20];
            mult_part_out06[318] <= P_10_5[28];
            mult_part_out06[319] <= P_3_10[28];
            mult_part_out06[320] <= P_11_5[13];
            mult_part_out06[321] <= P_11_4[38];
            mult_part_out06[322] <= P_11_5[15];
            mult_part_out06[323] <= P_4_10[15];
            mult_part_out06[324] <= P_11_5[17];
            mult_part_out06[325] <= P_15_2[22];
            mult_part_out06[326] <= P_11_5[19];
            mult_part_out06[327] <= P_5_10[2];
            mult_part_out06[328] <= P_10_6[14];
            mult_part_out06[329] <= P_10_5[39];
            mult_part_out06[330] <= P_8_7[26];
            mult_part_out06[331] <= P_9_7[10];
            mult_part_out06[332] <= P_4_10[24];
            mult_part_out06[333] <= P_8_8[5];
            mult_part_out06[334] <= P_12_5[10];
            mult_part_out06[335] <= P_7_9[0];
            mult_part_out06[336] <= P_12_4[36];
            mult_part_out06[337] <= P_14_4[3];
            mult_part_out06[338] <= P_14_4[4];
            mult_part_out06[339] <= P_12_5[15];
            mult_part_out06[340] <= P_13_4[23];
            mult_part_out06[341] <= P_7_8[30];
            mult_part_out06[342] <= P_6_9[24];
            mult_part_out06[343] <= P_8_8[15];
            mult_part_out06[344] <= P_7_9[9];
            mult_part_out06[345] <= P_5_10[20];
            mult_part_out06[346] <= P_9_8[1];
            mult_part_out06[347] <= P_14_4[13];
            mult_part_out06[348] <= P_9_8[3];
            mult_part_out06[349] <= P_6_9[31];
            mult_part_out06[350] <= P_8_8[22];
            mult_part_out06[351] <= P_5_10[26];
            mult_part_out06[352] <= P_12_5[28];
            mult_part_out06[353] <= P_15_4[2];
            mult_part_out06[354] <= P_9_8[9];
            mult_part_out06[355] <= P_6_9[37];
            mult_part_out06[356] <= P_9_8[11];
            mult_part_out06[357] <= P_8_8[29];
            mult_part_out06[358] <= P_14_4[24];
            mult_part_out06[359] <= P_14_5[1];
            mult_part_out06[360] <= P_7_10[1];
            mult_part_out06[361] <= P_14_4[27];
            mult_part_out06[362] <= P_12_5[38];
            mult_part_out06[363] <= P_11_6[32];
            mult_part_out06[364] <= P_6_10[22];
            mult_part_out06[365] <= P_13_5[24];
            mult_part_out06[366] <= P_13_6[1];
            mult_part_out06[367] <= P_7_9[32];
            mult_part_out06[368] <= P_8_8[40];
            mult_part_out06[369] <= P_9_9[0];
            mult_part_out06[370] <= P_12_6[22];
            mult_part_out06[371] <= P_12_6[23];
            mult_part_out06[372] <= P_12_6[24];
            mult_part_out06[373] <= P_14_5[15];
            mult_part_out06[374] <= P_15_4[23];
            mult_part_out06[375] <= P_12_7[3];
            mult_part_out06[376] <= P_9_8[31];
            mult_part_out06[377] <= P_8_10[1];
            mult_part_out06[378] <= P_9_9[9];
            mult_part_out06[379] <= P_12_6[31];
            mult_part_out06[380] <= P_12_6[32];
            mult_part_out06[381] <= P_15_5[6];
            mult_part_out06[382] <= P_13_6[17];
            mult_part_out06[383] <= P_12_6[35];
            mult_part_out06[384] <= P_9_8[39];
            mult_part_out06[385] <= P_10_8[23];
            mult_part_out06[386] <= P_15_5[11];
            mult_part_out06[387] <= P_11_8[8];
            mult_part_out06[388] <= P_7_10[29];
            mult_part_out06[389] <= P_15_5[14];
            mult_part_out06[390] <= P_11_7[35];
            mult_part_out06[391] <= P_13_7[2];
            mult_part_out06[392] <= P_12_7[20];
            mult_part_out06[393] <= P_10_9[7];
            mult_part_out06[394] <= P_14_5[36];
            mult_part_out06[395] <= P_13_7[6];
            mult_part_out06[396] <= P_11_8[17];
            mult_part_out06[397] <= P_14_6[15];
            mult_part_out06[398] <= P_14_5[40];
            mult_part_out06[399] <= P_11_8[20];
            mult_part_out06[400] <= P_12_8[4];
            mult_part_out06[401] <= P_14_6[19];
            mult_part_out06[402] <= P_12_8[6];
            mult_part_out06[403] <= P_13_6[38];
            mult_part_out06[404] <= P_10_9[18];
            mult_part_out06[405] <= P_12_7[33];
            mult_part_out06[406] <= P_10_9[20];
            mult_part_out06[407] <= P_11_9[4];
            mult_part_out06[408] <= P_10_9[22];
            mult_part_out06[409] <= P_9_10[16];
            mult_part_out06[410] <= P_14_7[4];
            mult_part_out06[411] <= P_13_7[22];
            mult_part_out06[412] <= P_12_8[16];
            mult_part_out06[413] <= P_12_8[17];
            mult_part_out06[414] <= P_12_8[18];
            mult_part_out06[415] <= P_12_8[19];
            mult_part_out06[416] <= P_11_9[13];
            mult_part_out06[417] <= P_14_7[11];
            mult_part_out06[418] <= P_11_8[39];
            mult_part_out06[419] <= P_13_7[30];
            mult_part_out06[420] <= P_15_6[21];
            mult_part_out06[421] <= P_14_7[15];
            mult_part_out06[422] <= P_12_8[26];
            mult_part_out06[423] <= P_11_9[20];
            mult_part_out06[424] <= P_13_8[11];
            mult_part_out06[425] <= P_13_7[36];
            mult_part_out06[426] <= P_11_9[23];
            mult_part_out06[427] <= P_12_8[31];
            mult_part_out06[428] <= P_11_10[1];
            mult_part_out06[429] <= P_15_7[6];
            mult_part_out06[430] <= P_10_10[20];
            mult_part_out06[431] <= P_12_9[11];
            mult_part_out06[432] <= P_13_8[19];
            mult_part_out06[433] <= P_12_8[37];
            mult_part_out06[434] <= P_11_10[7];
            mult_part_out06[435] <= P_15_7[12];
            mult_part_out06[436] <= P_15_7[13];
            mult_part_out06[437] <= P_14_8[7];
            mult_part_out06[438] <= P_13_9[1];
            mult_part_out06[439] <= P_11_10[12];
            mult_part_out06[440] <= P_12_9[20];
            mult_part_out06[441] <= P_13_9[4];
            mult_part_out06[442] <= P_13_8[29];
            mult_part_out06[443] <= P_13_9[6];
            mult_part_out06[444] <= P_13_9[7];
            mult_part_out06[445] <= P_14_7[39];
            mult_part_out06[446] <= P_12_9[26];
            mult_part_out06[447] <= P_12_10[3];
            mult_part_out06[448] <= P_15_8[1];
            mult_part_out06[449] <= P_12_10[5];
            mult_part_out06[450] <= P_15_8[3];
            mult_part_out06[451] <= P_11_10[24];
            mult_part_out06[452] <= P_12_10[8];
            mult_part_out06[453] <= P_13_8[40];
            mult_part_out06[454] <= P_14_9[0];
            mult_part_out06[455] <= P_15_8[8];
            mult_part_out06[456] <= P_13_9[19];
            mult_part_out06[457] <= P_12_10[13];
            mult_part_out06[458] <= P_12_9[38];
            mult_part_out06[459] <= P_12_9[39];

            mult_part_out07[72] <= P_0_3[0];
            mult_part_out07[73] <= P_1_2[8];
            mult_part_out07[74] <= P_0_2[26];
            mult_part_out07[75] <= P_3_0[24];
            mult_part_out07[76] <= P_0_2[28];
            mult_part_out07[77] <= P_0_3[5];
            mult_part_out07[78] <= P_0_3[6];
            mult_part_out07[79] <= P_3_1[4];
            mult_part_out07[80] <= P_2_1[22];
            mult_part_out07[81] <= P_1_2[16];
            mult_part_out07[82] <= P_3_0[31];
            mult_part_out07[83] <= P_3_1[8];
            mult_part_out07[84] <= P_4_0[16];
            mult_part_out07[85] <= P_2_1[27];
            mult_part_out07[86] <= P_5_0[1];
            mult_part_out07[87] <= P_2_2[5];
            mult_part_out07[88] <= P_1_2[23];
            mult_part_out07[89] <= P_5_0[4];
            mult_part_out07[90] <= P_1_3[1];
            mult_part_out07[91] <= P_1_3[2];
            mult_part_out07[92] <= P_2_2[10];
            mult_part_out07[93] <= P_3_1[18];
            mult_part_out07[94] <= P_0_3[22];
            mult_part_out07[95] <= P_5_0[10];
            mult_part_out07[96] <= P_2_2[14];
            mult_part_out07[97] <= P_1_3[8];
            mult_part_out07[98] <= P_4_1[6];
            mult_part_out07[99] <= P_0_3[27];
            mult_part_out07[100] <= P_4_1[8];
            mult_part_out07[101] <= P_1_2[36];
            mult_part_out07[102] <= P_1_2[37];
            mult_part_out07[103] <= P_4_0[35];
            mult_part_out07[104] <= P_2_2[22];
            mult_part_out07[105] <= P_0_4[9];
            mult_part_out07[106] <= P_0_4[10];
            mult_part_out07[107] <= P_0_3[35];
            mult_part_out07[108] <= P_4_0[40];
            mult_part_out07[109] <= P_0_3[37];
            mult_part_out07[110] <= P_2_2[28];
            mult_part_out07[111] <= P_0_3[39];
            mult_part_out07[112] <= P_0_4[16];
            mult_part_out07[113] <= P_3_1[38];
            mult_part_out07[114] <= P_5_1[5];
            mult_part_out07[115] <= P_5_1[6];
            mult_part_out07[116] <= P_4_1[24];
            mult_part_out07[117] <= P_2_3[11];
            mult_part_out07[118] <= P_1_3[29];
            mult_part_out07[119] <= P_2_3[13];
            mult_part_out07[120] <= P_5_1[11];
            mult_part_out07[121] <= P_5_0[36];
            mult_part_out07[122] <= P_3_2[23];
            mult_part_out07[123] <= P_2_3[17];
            mult_part_out07[124] <= P_6_0[22];
            mult_part_out07[125] <= P_1_4[12];
            mult_part_out07[126] <= P_5_1[17];
            mult_part_out07[127] <= P_1_4[14];
            mult_part_out07[128] <= P_0_4[32];
            mult_part_out07[129] <= P_6_1[3];
            mult_part_out07[130] <= P_7_0[11];
            mult_part_out07[131] <= P_2_3[25];
            mult_part_out07[132] <= P_5_1[23];
            mult_part_out07[133] <= P_5_2[0];
            mult_part_out07[134] <= P_7_0[15];
            mult_part_out07[135] <= P_3_3[12];
            mult_part_out07[136] <= P_8_0[0];
            mult_part_out07[137] <= P_5_2[4];
            mult_part_out07[138] <= P_3_3[15];
            mult_part_out07[139] <= P_8_0[3];
            mult_part_out07[140] <= P_1_5[3];
            mult_part_out07[141] <= P_2_3[35];
            mult_part_out07[142] <= P_6_1[16];
            mult_part_out07[143] <= P_2_4[13];
            mult_part_out07[144] <= P_4_3[4];
            mult_part_out07[145] <= P_0_6[1];
            mult_part_out07[146] <= P_5_1[37];
            mult_part_out07[147] <= P_0_5[27];
            mult_part_out07[148] <= P_1_5[11];
            mult_part_out07[149] <= P_6_1[23];
            mult_part_out07[150] <= P_7_1[7];
            mult_part_out07[151] <= P_7_0[32];
            mult_part_out07[152] <= P_1_4[39];
            mult_part_out07[153] <= P_8_0[17];
            mult_part_out07[154] <= P_2_4[24];
            mult_part_out07[155] <= P_2_4[25];
            mult_part_out07[156] <= P_3_3[33];
            mult_part_out07[157] <= P_7_1[14];
            mult_part_out07[158] <= P_3_3[35];
            mult_part_out07[159] <= P_2_5[5];
            mult_part_out07[160] <= P_6_2[10];
            mult_part_out07[161] <= P_1_6[0];
            mult_part_out07[162] <= P_3_4[15];
            mult_part_out07[163] <= P_1_6[2];
            mult_part_out07[164] <= P_7_1[21];
            mult_part_out07[165] <= P_8_1[5];
            mult_part_out07[166] <= P_0_6[22];
            mult_part_out07[167] <= P_3_4[20];
            mult_part_out07[168] <= P_8_0[32];
            mult_part_out07[169] <= P_4_3[29];
            mult_part_out07[170] <= P_1_6[9];
            mult_part_out07[171] <= P_2_5[17];
            mult_part_out07[172] <= P_5_3[15];
            mult_part_out07[173] <= P_0_6[29];
            mult_part_out07[174] <= P_0_6[30];
            mult_part_out07[175] <= P_6_3[1];
            mult_part_out07[176] <= P_1_6[15];
            mult_part_out07[177] <= P_10_0[7];
            mult_part_out07[178] <= P_0_6[34];
            mult_part_out07[179] <= P_2_6[1];
            mult_part_out07[180] <= P_1_6[19];
            mult_part_out07[181] <= P_9_0[28];
            mult_part_out07[182] <= P_0_6[38];
            mult_part_out07[183] <= P_0_7[15];
            mult_part_out07[184] <= P_4_4[20];
            mult_part_out07[185] <= P_3_5[14];
            mult_part_out07[186] <= P_3_4[39];
            mult_part_out07[187] <= P_9_1[10];
            mult_part_out07[188] <= P_11_0[1];
            mult_part_out07[189] <= P_8_2[5];
            mult_part_out07[190] <= P_2_5[36];
            mult_part_out07[191] <= P_5_4[10];
            mult_part_out07[192] <= P_5_4[11];
            mult_part_out07[193] <= P_10_0[23];
            mult_part_out07[194] <= P_8_1[34];
            mult_part_out07[195] <= P_3_6[0];
            mult_part_out07[196] <= P_11_0[9];
            mult_part_out07[197] <= P_2_6[19];
            mult_part_out07[198] <= P_1_6[37];
            mult_part_out07[199] <= P_0_8[7];
            mult_part_out07[200] <= P_7_3[9];
            mult_part_out07[201] <= P_6_3[27];
            mult_part_out07[202] <= P_3_5[31];
            mult_part_out07[203] <= P_10_1[9];
            mult_part_out07[204] <= P_2_7[2];
            mult_part_out07[205] <= P_6_3[31];
            mult_part_out07[206] <= P_6_3[32];
            mult_part_out07[207] <= P_2_7[5];
            mult_part_out07[208] <= P_3_6[13];
            mult_part_out07[209] <= P_5_4[28];
            mult_part_out07[210] <= P_5_4[29];
            mult_part_out07[211] <= P_2_7[9];
            mult_part_out07[212] <= P_2_7[10];
            mult_part_out07[213] <= P_0_8[21];
            mult_part_out07[214] <= P_6_3[40];
            mult_part_out07[215] <= P_4_6[3];
            mult_part_out07[216] <= P_5_5[11];
            mult_part_out07[217] <= P_11_0[30];
            mult_part_out07[218] <= P_12_0[14];
            mult_part_out07[219] <= P_3_7[0];
            mult_part_out07[220] <= P_4_5[32];
            mult_part_out07[221] <= P_10_2[3];
            mult_part_out07[222] <= P_6_4[24];
            mult_part_out07[223] <= P_0_8[31];
            mult_part_out07[224] <= P_11_1[13];
            mult_part_out07[225] <= P_6_4[27];
            mult_part_out07[226] <= P_0_9[10];
            mult_part_out07[227] <= P_13_0[6];
            mult_part_out07[228] <= P_4_5[40];
            mult_part_out07[229] <= P_12_0[25];
            mult_part_out07[230] <= P_1_8[21];
            mult_part_out07[231] <= P_2_7[29];
            mult_part_out07[232] <= P_2_7[30];
            mult_part_out07[233] <= P_1_8[24];
            mult_part_out07[234] <= P_0_9[18];
            mult_part_out07[235] <= P_7_4[20];
            mult_part_out07[236] <= P_1_8[27];
            mult_part_out07[237] <= P_8_4[5];
            mult_part_out07[238] <= P_8_3[30];
            mult_part_out07[239] <= P_4_7[3];
            mult_part_out07[240] <= P_12_1[12];
            mult_part_out07[241] <= P_7_4[26];
            mult_part_out07[242] <= P_13_0[21];
            mult_part_out07[243] <= P_0_10[3];
            mult_part_out07[244] <= P_6_5[22];
            mult_part_out07[245] <= P_3_7[26];
            mult_part_out07[246] <= P_6_6[0];
            mult_part_out07[247] <= P_7_5[8];
            mult_part_out07[248] <= P_1_9[15];
            mult_part_out07[249] <= P_11_2[14];
            mult_part_out07[250] <= P_4_6[38];
            mult_part_out07[251] <= P_12_1[23];
            mult_part_out07[252] <= P_0_9[36];
            mult_part_out07[253] <= P_4_7[17];
            mult_part_out07[254] <= P_3_7[35];
            mult_part_out07[255] <= P_0_10[15];
            mult_part_out07[256] <= P_14_0[18];
            mult_part_out07[257] <= P_13_0[36];
            mult_part_out07[258] <= P_12_2[6];
            mult_part_out07[259] <= P_12_1[31];
            mult_part_out07[260] <= P_1_10[3];
            mult_part_out07[261] <= P_13_0[40];
            mult_part_out07[262] <= P_5_6[33];
            mult_part_out07[263] <= P_7_6[0];
            mult_part_out07[264] <= P_5_6[35];
            mult_part_out07[265] <= P_4_7[29];
            mult_part_out07[266] <= P_12_1[38];
            mult_part_out07[267] <= P_7_5[28];
            mult_part_out07[268] <= P_12_2[16];
            mult_part_out07[269] <= P_1_10[12];
            mult_part_out07[270] <= P_8_5[14];
            mult_part_out07[271] <= P_11_3[12];
            mult_part_out07[272] <= P_13_2[3];
            mult_part_out07[273] <= P_7_5[34];
            mult_part_out07[274] <= P_11_2[39];
            mult_part_out07[275] <= P_3_9[8];
            mult_part_out07[276] <= P_14_1[14];
            mult_part_out07[277] <= P_7_6[14];
            mult_part_out07[278] <= P_7_6[15];
            mult_part_out07[279] <= P_5_7[26];
            mult_part_out07[280] <= P_13_1[35];
            mult_part_out07[281] <= P_11_3[22];
            mult_part_out07[282] <= P_8_6[2];
            mult_part_out07[283] <= P_4_8[23];
            mult_part_out07[284] <= P_11_3[25];
            mult_part_out07[285] <= P_12_2[33];
            mult_part_out07[286] <= P_15_1[7];
            mult_part_out07[287] <= P_14_2[1];
            mult_part_out07[288] <= P_8_5[32];
            mult_part_out07[289] <= P_9_5[16];
            mult_part_out07[290] <= P_9_5[17];
            mult_part_out07[291] <= P_9_5[18];
            mult_part_out07[292] <= P_3_9[25];
            mult_part_out07[293] <= P_11_3[34];
            mult_part_out07[294] <= P_11_3[35];
            mult_part_out07[295] <= P_3_9[28];
            mult_part_out07[296] <= P_5_8[19];
            mult_part_out07[297] <= P_4_9[13];
            mult_part_out07[298] <= P_13_2[29];
            mult_part_out07[299] <= P_11_3[40];
            mult_part_out07[300] <= P_14_1[38];
            mult_part_out07[301] <= P_13_3[8];
            mult_part_out07[302] <= P_3_10[11];
            mult_part_out07[303] <= P_6_8[9];
            mult_part_out07[304] <= P_13_3[11];
            mult_part_out07[305] <= P_11_4[22];
            mult_part_out07[306] <= P_8_7[2];
            mult_part_out07[307] <= P_4_9[23];
            mult_part_out07[308] <= P_13_2[39];
            mult_part_out07[309] <= P_8_7[5];
            mult_part_out07[310] <= P_6_7[40];
            mult_part_out07[311] <= P_12_4[11];
            mult_part_out07[312] <= P_12_3[36];
            mult_part_out07[313] <= P_12_4[13];
            mult_part_out07[314] <= P_14_3[4];
            mult_part_out07[315] <= P_3_10[24];
            mult_part_out07[316] <= P_12_4[16];
            mult_part_out07[317] <= P_10_5[27];
            mult_part_out07[318] <= P_9_6[21];
            mult_part_out07[319] <= P_4_10[11];
            mult_part_out07[320] <= P_14_2[34];
            mult_part_out07[321] <= P_12_4[21];
            mult_part_out07[322] <= P_6_9[4];
            mult_part_out07[323] <= P_3_10[32];
            mult_part_out07[324] <= P_13_4[7];
            mult_part_out07[325] <= P_6_8[31];
            mult_part_out07[326] <= P_12_4[26];
            mult_part_out07[327] <= P_5_9[26];
            mult_part_out07[328] <= P_5_10[3];
            mult_part_out07[329] <= P_15_3[2];
            mult_part_out07[330] <= P_8_8[2];
            mult_part_out07[331] <= P_11_5[24];
            mult_part_out07[332] <= P_6_8[38];
            mult_part_out07[333] <= P_12_4[33];
            mult_part_out07[334] <= P_8_7[30];
            mult_part_out07[335] <= P_8_8[7];
            mult_part_out07[336] <= P_14_3[26];
            mult_part_out07[337] <= P_8_7[33];
            mult_part_out07[338] <= P_6_9[20];
            mult_part_out07[339] <= P_12_4[39];
            mult_part_out07[340] <= P_11_5[33];
            mult_part_out07[341] <= P_9_7[20];
            mult_part_out07[342] <= P_14_4[8];
            mult_part_out07[343] <= P_6_9[25];
            mult_part_out07[344] <= P_6_9[26];
            mult_part_out07[345] <= P_6_10[3];
            mult_part_out07[346] <= P_12_5[22];
            mult_part_out07[347] <= P_6_10[5];
            mult_part_out07[348] <= P_9_7[27];
            mult_part_out07[349] <= P_7_8[38];
            mult_part_out07[350] <= P_5_10[25];
            mult_part_out07[351] <= P_7_9[16];
            mult_part_out07[352] <= P_9_7[31];
            mult_part_out07[353] <= P_7_9[18];
            mult_part_out07[354] <= P_8_9[2];
            mult_part_out07[355] <= P_9_8[10];
            mult_part_out07[356] <= P_13_5[15];
            mult_part_out07[357] <= P_9_7[36];
            mult_part_out07[358] <= P_9_7[37];
            mult_part_out07[359] <= P_9_8[14];
            mult_part_out07[360] <= P_6_10[18];
            mult_part_out07[361] <= P_7_9[26];
            mult_part_out07[362] <= P_13_5[21];
            mult_part_out07[363] <= P_14_4[29];
            mult_part_out07[364] <= P_10_7[26];
            mult_part_out07[365] <= P_13_6[0];
            mult_part_out07[366] <= P_9_8[21];
            mult_part_out07[367] <= P_8_8[39];
            mult_part_out07[368] <= P_7_10[9];
            mult_part_out07[369] <= P_6_10[27];
            mult_part_out07[370] <= P_7_10[11];
            mult_part_out07[371] <= P_13_6[6];
            mult_part_out07[372] <= P_15_4[21];
            mult_part_out07[373] <= P_14_4[39];
            mult_part_out07[374] <= P_7_10[15];
            mult_part_out07[375] <= P_9_9[6];
            mult_part_out07[376] <= P_15_5[1];
            mult_part_out07[377] <= P_7_10[18];
            mult_part_out07[378] <= P_7_10[19];
            mult_part_out07[379] <= P_15_5[4];
            mult_part_out07[380] <= P_7_10[21];
            mult_part_out07[381] <= P_11_8[2];
            mult_part_out07[382] <= P_12_6[34];
            mult_part_out07[383] <= P_8_9[31];
            mult_part_out07[384] <= P_12_6[36];
            mult_part_out07[385] <= P_8_10[9];
            mult_part_out07[386] <= P_7_10[27];
            mult_part_out07[387] <= P_7_10[28];
            mult_part_out07[388] <= P_11_8[9];
            mult_part_out07[389] <= P_11_8[10];
            mult_part_out07[390] <= P_15_5[15];
            mult_part_out07[391] <= P_14_5[33];
            mult_part_out07[392] <= P_11_7[37];
            mult_part_out07[393] <= P_8_10[17];
            mult_part_out07[394] <= P_9_9[25];
            mult_part_out07[395] <= P_8_10[19];
            mult_part_out07[396] <= P_14_5[38];
            mult_part_out07[397] <= P_10_8[35];
            mult_part_out07[398] <= P_15_5[23];
            mult_part_out07[399] <= P_13_7[10];
            mult_part_out07[400] <= P_10_8[38];
            mult_part_out07[401] <= P_10_8[39];
            mult_part_out07[402] <= P_15_6[3];
            mult_part_out07[403] <= P_11_9[0];
            mult_part_out07[404] <= P_9_10[11];
            mult_part_out07[405] <= P_12_8[9];
            mult_part_out07[406] <= P_13_7[17];
            mult_part_out07[407] <= P_11_8[28];
            mult_part_out07[408] <= P_15_6[9];
            mult_part_out07[409] <= P_12_8[13];
            mult_part_out07[410] <= P_15_6[11];
            mult_part_out07[411] <= P_12_8[15];
            mult_part_out07[412] <= P_14_7[6];
            mult_part_out07[413] <= P_13_8[0];
            mult_part_out07[414] <= P_9_10[21];
            mult_part_out07[415] <= P_13_8[2];
            mult_part_out07[416] <= P_12_8[20];
            mult_part_out07[417] <= P_10_9[31];
            mult_part_out07[418] <= P_15_6[19];
            mult_part_out07[419] <= P_10_9[33];
            mult_part_out07[420] <= P_13_7[31];
            mult_part_out07[421] <= P_15_6[22];
            mult_part_out07[422] <= P_11_9[19];
            mult_part_out07[423] <= P_12_8[27];
            mult_part_out07[424] <= P_14_7[18];
            mult_part_out07[425] <= P_12_8[29];
            mult_part_out07[426] <= P_12_8[30];
            mult_part_out07[427] <= P_12_9[7];
            mult_part_out07[428] <= P_15_7[5];
            mult_part_out07[429] <= P_11_10[2];
            mult_part_out07[430] <= P_12_8[34];
            mult_part_out07[431] <= P_10_10[21];
            mult_part_out07[432] <= P_12_9[12];
            mult_part_out07[433] <= P_14_8[3];
            mult_part_out07[434] <= P_12_9[14];
            mult_part_out07[435] <= P_14_7[29];
            mult_part_out07[436] <= P_14_7[30];
            mult_part_out07[437] <= P_10_10[27];
            mult_part_out07[438] <= P_14_7[32];
            mult_part_out07[439] <= P_10_10[29];
            mult_part_out07[440] <= P_11_10[13];
            mult_part_out07[441] <= P_11_10[14];
            mult_part_out07[442] <= P_12_9[22];
            mult_part_out07[443] <= P_11_9[40];
            mult_part_out07[444] <= P_14_8[14];
            mult_part_out07[445] <= P_12_10[1];
            mult_part_out07[446] <= P_12_10[2];
            mult_part_out07[447] <= P_13_8[34];

            mult_part_out08[85] <= P_3_0[34];
            mult_part_out08[86] <= P_4_0[18];
            mult_part_out08[87] <= P_3_0[36];
            mult_part_out08[88] <= P_2_2[6];
            mult_part_out08[89] <= P_3_0[38];
            mult_part_out08[90] <= P_3_0[39];
            mult_part_out08[91] <= P_2_2[9];
            mult_part_out08[92] <= P_4_1[0];
            mult_part_out08[93] <= P_1_2[28];
            mult_part_out08[94] <= P_4_1[2];
            mult_part_out08[95] <= P_3_1[20];
            mult_part_out08[96] <= P_1_2[31];
            mult_part_out08[97] <= P_4_1[5];
            mult_part_out08[98] <= P_1_3[9];
            mult_part_out08[99] <= P_4_1[7];
            mult_part_out08[100] <= P_1_2[35];
            mult_part_out08[101] <= P_0_4[5];
            mult_part_out08[102] <= P_3_2[3];
            mult_part_out08[103] <= P_2_2[21];
            mult_part_out08[104] <= P_0_4[8];
            mult_part_out08[105] <= P_1_2[40];
            mult_part_out08[106] <= P_3_2[7];
            mult_part_out08[107] <= P_0_4[11];
            mult_part_out08[108] <= P_0_4[12];
            mult_part_out08[109] <= P_3_1[34];
            mult_part_out08[110] <= P_0_3[38];
            mult_part_out08[111] <= P_1_3[22];
            mult_part_out08[112] <= P_4_1[20];
            mult_part_out08[113] <= P_0_4[17];
            mult_part_out08[114] <= P_2_3[8];
            mult_part_out08[115] <= P_4_1[23];
            mult_part_out08[116] <= P_4_2[0];
            mult_part_out08[117] <= P_4_2[1];
            mult_part_out08[118] <= P_0_4[22];
            mult_part_out08[119] <= P_5_1[10];
            mult_part_out08[120] <= P_5_0[35];
            mult_part_out08[121] <= P_1_3[32];
            mult_part_out08[122] <= P_0_5[2];
            mult_part_out08[123] <= P_4_2[7];
            mult_part_out08[124] <= P_1_3[35];
            mult_part_out08[125] <= P_3_2[26];
            mult_part_out08[126] <= P_6_1[0];
            mult_part_out08[127] <= P_2_3[21];
            mult_part_out08[128] <= P_6_1[2];
            mult_part_out08[129] <= P_6_0[27];
            mult_part_out08[130] <= P_4_1[38];
            mult_part_out08[131] <= P_2_4[1];
            mult_part_out08[132] <= P_3_3[9];
            mult_part_out08[133] <= P_2_3[27];
            mult_part_out08[134] <= P_2_3[28];
            mult_part_out08[135] <= P_0_4[39];
            mult_part_out08[136] <= P_3_3[13];
            mult_part_out08[137] <= P_0_5[17];
            mult_part_out08[138] <= P_6_0[36];
            mult_part_out08[139] <= P_1_4[26];
            mult_part_out08[140] <= P_4_2[24];
            mult_part_out08[141] <= P_2_4[11];
            mult_part_out08[142] <= P_4_3[2];
            mult_part_out08[143] <= P_0_5[23];
            mult_part_out08[144] <= P_5_1[35];
            mult_part_out08[145] <= P_4_2[29];
            mult_part_out08[146] <= P_6_1[20];
            mult_part_out08[147] <= P_7_1[4];
            mult_part_out08[148] <= P_5_1[39];
            mult_part_out08[149] <= P_5_1[40];
            mult_part_out08[150] <= P_8_0[14];
            mult_part_out08[151] <= P_8_0[15];
            mult_part_out08[152] <= P_4_3[12];
            mult_part_out08[153] <= P_4_3[13];
            mult_part_out08[154] <= P_0_5[34];
            mult_part_out08[155] <= P_7_0[36];
            mult_part_out08[156] <= P_5_2[23];
            mult_part_out08[157] <= P_6_1[31];
            mult_part_out08[158] <= P_8_0[22];
            mult_part_out08[159] <= P_3_3[36];
            mult_part_out08[160] <= P_3_4[13];
            mult_part_out08[161] <= P_5_3[4];
            mult_part_out08[162] <= P_6_1[36];
            mult_part_out08[163] <= P_4_3[23];
            mult_part_out08[164] <= P_9_0[11];
            mult_part_out08[165] <= P_4_4[1];
            mult_part_out08[166] <= P_6_2[16];
            mult_part_out08[167] <= P_4_4[3];
            mult_part_out08[168] <= P_7_2[1];
            mult_part_out08[169] <= P_8_0[33];
            mult_part_out08[170] <= P_2_5[16];
            mult_part_out08[171] <= P_5_3[14];
            mult_part_out08[172] <= P_4_4[8];
            mult_part_out08[173] <= P_10_0[3];
            mult_part_out08[174] <= P_1_6[13];
            mult_part_out08[175] <= P_0_7[7];
            mult_part_out08[176] <= P_2_5[22];
            mult_part_out08[177] <= P_7_1[34];
            mult_part_out08[178] <= P_3_4[31];
            mult_part_out08[179] <= P_6_2[29];
            mult_part_out08[180] <= P_8_1[20];
            mult_part_out08[181] <= P_10_0[11];
            mult_part_out08[182] <= P_0_7[14];
            mult_part_out08[183] <= P_9_0[30];
            mult_part_out08[184] <= P_10_0[14];
            mult_part_out08[185] <= P_10_0[15];
            mult_part_out08[186] <= P_5_3[29];
            mult_part_out08[187] <= P_5_4[6];
            mult_part_out08[188] <= P_9_0[35];
            mult_part_out08[189] <= P_11_0[2];
            mult_part_out08[190] <= P_11_0[3];
            mult_part_out08[191] <= P_11_0[4];
            mult_part_out08[192] <= P_1_7[7];
            mult_part_out08[193] <= P_9_0[40];
            mult_part_out08[194] <= P_10_0[24];
            mult_part_out08[195] <= P_5_4[14];
            mult_part_out08[196] <= P_4_5[8];
            mult_part_out08[197] <= P_6_3[23];
            mult_part_out08[198] <= P_11_0[11];
            mult_part_out08[199] <= P_6_4[1];
            mult_part_out08[200] <= P_2_6[22];
            mult_part_out08[201] <= P_9_2[0];
            mult_part_out08[202] <= P_10_1[8];
            mult_part_out08[203] <= P_1_7[18];
            mult_part_out08[204] <= P_3_6[9];
            mult_part_out08[205] <= P_11_0[18];
            mult_part_out08[206] <= P_11_0[19];
            mult_part_out08[207] <= P_8_2[23];
            mult_part_out08[208] <= P_9_2[7];
            mult_part_out08[209] <= P_2_7[7];
            mult_part_out08[210] <= P_8_3[2];
            mult_part_out08[211] <= P_8_3[3];
            mult_part_out08[212] <= P_1_8[3];
            mult_part_out08[213] <= P_1_8[4];
            mult_part_out08[214] <= P_4_5[26];
            mult_part_out08[215] <= P_2_7[13];
            mult_part_out08[216] <= P_2_7[14];
            mult_part_out08[217] <= P_6_4[19];
            mult_part_out08[218] <= P_8_3[10];
            mult_part_out08[219] <= P_11_1[8];
            mult_part_out08[220] <= P_11_0[33];
            mult_part_out08[221] <= P_12_0[17];
            mult_part_out08[222] <= P_3_6[27];
            mult_part_out08[223] <= P_13_0[2];
            mult_part_out08[224] <= P_11_0[37];
            mult_part_out08[225] <= P_1_8[16];
            mult_part_out08[226] <= P_6_4[28];
            mult_part_out08[227] <= P_6_5[5];
            mult_part_out08[228] <= P_2_8[2];
            mult_part_out08[229] <= P_12_1[1];
            mult_part_out08[230] <= P_3_7[11];
            mult_part_out08[231] <= P_3_6[36];
            mult_part_out08[232] <= P_1_8[23];
            mult_part_out08[233] <= P_0_9[17];
            mult_part_out08[234] <= P_6_5[12];
            mult_part_out08[235] <= P_12_0[31];
            mult_part_out08[236] <= P_9_2[35];
            mult_part_out08[237] <= P_2_7[35];
            mult_part_out08[238] <= P_2_8[12];
            mult_part_out08[239] <= P_10_2[21];
            mult_part_out08[240] <= P_9_3[15];
            mult_part_out08[241] <= P_0_9[25];
            mult_part_out08[242] <= P_7_4[27];
            mult_part_out08[243] <= P_13_0[22];
            mult_part_out08[244] <= P_3_7[25];
            mult_part_out08[245] <= P_2_8[19];
            mult_part_out08[246] <= P_0_10[6];
            mult_part_out08[247] <= P_11_2[12];
            mult_part_out08[248] <= P_2_8[22];
            mult_part_out08[249] <= P_13_1[4];
            mult_part_out08[250] <= P_13_1[5];
            mult_part_out08[251] <= P_10_3[9];
            mult_part_out08[252] <= P_3_8[9];
            mult_part_out08[253] <= P_5_6[24];
            mult_part_out08[254] <= P_10_2[36];
            mult_part_out08[255] <= P_13_0[34];
            mult_part_out08[256] <= P_3_8[13];
            mult_part_out08[257] <= P_15_0[2];
            mult_part_out08[258] <= P_2_8[32];
            mult_part_out08[259] <= P_13_0[38];
            mult_part_out08[260] <= P_5_6[31];
            mult_part_out08[261] <= P_9_4[12];
            mult_part_out08[262] <= P_8_5[6];
            mult_part_out08[263] <= P_9_4[14];
            mult_part_out08[264] <= P_6_6[18];
            mult_part_out08[265] <= P_8_4[33];
            mult_part_out08[266] <= P_4_7[30];
            mult_part_out08[267] <= P_14_0[29];
            mult_part_out08[268] <= P_2_9[18];
            mult_part_out08[269] <= P_14_0[31];
            mult_part_out08[270] <= P_14_0[32];
            mult_part_out08[271] <= P_6_7[1];
            mult_part_out08[272] <= P_10_3[30];
            mult_part_out08[273] <= P_3_9[6];
            mult_part_out08[274] <= P_5_7[21];
            mult_part_out08[275] <= P_11_2[40];
            mult_part_out08[276] <= P_3_9[9];
            mult_part_out08[277] <= P_14_0[39];
            mult_part_out08[278] <= P_13_1[33];
            mult_part_out08[279] <= P_7_5[40];
            mult_part_out08[280] <= P_5_8[3];
            mult_part_out08[281] <= P_9_5[8];
            mult_part_out08[282] <= P_10_4[16];
            mult_part_out08[283] <= P_14_1[21];
            mult_part_out08[284] <= P_4_9[0];
            mult_part_out08[285] <= P_15_1[6];
            mult_part_out08[286] <= P_13_2[17];
            mult_part_out08[287] <= P_15_1[8];
            mult_part_out08[288] <= P_11_4[5];
            mult_part_out08[289] <= P_12_2[37];
            mult_part_out08[290] <= P_13_2[21];
            mult_part_out08[291] <= P_3_10[0];
            mult_part_out08[292] <= P_10_5[2];
            mult_part_out08[293] <= P_8_6[13];
            mult_part_out08[294] <= P_8_6[14];
            mult_part_out08[295] <= P_9_5[22];
            mult_part_out08[296] <= P_15_1[17];
            mult_part_out08[297] <= P_10_5[7];
            mult_part_out08[298] <= P_9_5[25];
            mult_part_out08[299] <= P_2_10[25];
            mult_part_out08[300] <= P_14_2[14];
            mult_part_out08[301] <= P_10_4[35];
            mult_part_out08[302] <= P_5_9[1];
            mult_part_out08[303] <= P_10_4[37];
            mult_part_out08[304] <= P_6_7[34];
            mult_part_out08[305] <= P_2_10[31];
            mult_part_out08[306] <= P_9_6[9];
            mult_part_out08[307] <= P_3_9[40];
            mult_part_out08[308] <= P_4_9[24];
            mult_part_out08[309] <= P_4_10[1];
            mult_part_out08[310] <= P_8_7[6];
            mult_part_out08[311] <= P_13_3[18];
            mult_part_out08[312] <= P_10_5[22];
            mult_part_out08[313] <= P_14_2[27];
            mult_part_out08[314] <= P_15_2[11];
            mult_part_out08[315] <= P_9_6[18];
            mult_part_out08[316] <= P_7_7[29];
            mult_part_out08[317] <= P_5_8[40];
            mult_part_out08[318] <= P_7_7[31];
            mult_part_out08[319] <= P_5_9[18];
            mult_part_out08[320] <= P_8_6[40];
            mult_part_out08[321] <= P_9_6[24];
            mult_part_out08[322] <= P_8_7[18];
            mult_part_out08[323] <= P_14_3[13];
            mult_part_out08[324] <= P_12_4[24];
            mult_part_out08[325] <= P_14_2[39];
            mult_part_out08[326] <= P_6_8[32];
            mult_part_out08[327] <= P_10_5[37];
            mult_part_out08[328] <= P_7_8[17];
            mult_part_out08[329] <= P_11_5[22];
            mult_part_out08[330] <= P_5_10[5];
            mult_part_out08[331] <= P_15_3[4];
            mult_part_out08[332] <= P_9_7[11];
            mult_part_out08[333] <= P_13_3[40];
            mult_part_out08[334] <= P_5_9[33];
            mult_part_out08[335] <= P_11_6[4];
            mult_part_out08[336] <= P_8_8[8];
            mult_part_out08[337] <= P_12_4[37];
            mult_part_out08[338] <= P_5_9[37];
            mult_part_out08[339] <= P_5_9[38];
            mult_part_out08[340] <= P_12_4[40];
            mult_part_out08[341] <= P_7_9[6];
            mult_part_out08[342] <= P_10_7[4];
            mult_part_out08[343] <= P_14_3[33];
            mult_part_out08[344] <= P_13_4[27];
            mult_part_out08[345] <= P_7_9[10];
            mult_part_out08[346] <= P_11_6[15];
            mult_part_out08[347] <= P_8_8[19];
            mult_part_out08[348] <= P_13_4[31];
            mult_part_out08[349] <= P_10_7[11];
            mult_part_out08[350] <= P_10_7[12];
            mult_part_out08[351] <= P_10_7[13];
            mult_part_out08[352] <= P_10_6[38];
            mult_part_out08[353] <= P_9_7[32];
            mult_part_out08[354] <= P_14_4[20];
            mult_part_out08[355] <= P_10_7[17];
            mult_part_out08[356] <= P_11_6[25];
            mult_part_out08[357] <= P_12_5[33];
            mult_part_out08[358] <= P_11_6[27];
            mult_part_out08[359] <= P_14_4[25];
            mult_part_out08[360] <= P_9_8[15];
            mult_part_out08[361] <= P_9_7[40];
            mult_part_out08[362] <= P_12_6[14];
            mult_part_out08[363] <= P_15_4[12];
            mult_part_out08[364] <= P_11_7[9];
            mult_part_out08[365] <= P_11_7[10];
            mult_part_out08[366] <= P_12_6[18];
            mult_part_out08[367] <= P_6_10[25];
            mult_part_out08[368] <= P_6_10[26];
            mult_part_out08[369] <= P_7_10[10];
            mult_part_out08[370] <= P_13_6[5];
            mult_part_out08[371] <= P_9_9[2];
            mult_part_out08[372] <= P_13_6[7];
            mult_part_out08[373] <= P_15_4[22];
            mult_part_out08[374] <= P_9_9[5];
            mult_part_out08[375] <= P_7_10[16];
            mult_part_out08[376] <= P_14_5[18];
            mult_part_out08[377] <= P_9_8[32];
            mult_part_out08[378] <= P_11_7[23];
            mult_part_out08[379] <= P_14_5[21];
            mult_part_out08[380] <= P_8_10[4];
            mult_part_out08[381] <= P_14_5[23];
            mult_part_out08[382] <= P_14_5[24];
            mult_part_out08[383] <= P_13_6[18];
            mult_part_out08[384] <= P_14_5[26];
            mult_part_out08[385] <= P_15_5[10];
            mult_part_out08[386] <= P_14_6[4];
            mult_part_out08[387] <= P_12_7[15];
            mult_part_out08[388] <= P_12_6[40];
            mult_part_out08[389] <= P_13_7[0];
            mult_part_out08[390] <= P_14_5[32];
            mult_part_out08[391] <= P_9_9[22];
            mult_part_out08[392] <= P_10_9[6];
            mult_part_out08[393] <= P_12_7[21];
            mult_part_out08[394] <= P_14_6[12];
            mult_part_out08[395] <= P_15_5[20];
            mult_part_out08[396] <= P_15_5[21];
            mult_part_out08[397] <= P_15_5[22];
            mult_part_out08[398] <= P_9_9[29];
            mult_part_out08[399] <= P_8_10[23];
            mult_part_out08[400] <= P_9_10[7];
            mult_part_out08[401] <= P_12_7[29];
            mult_part_out08[402] <= P_9_10[9];
            mult_part_out08[403] <= P_8_10[27];
            mult_part_out08[404] <= P_15_6[5];
            mult_part_out08[405] <= P_14_6[23];
            mult_part_out08[406] <= P_9_9[37];
            mult_part_out08[407] <= P_12_7[35];
            mult_part_out08[408] <= P_11_8[29];
            mult_part_out08[409] <= P_11_9[6];
            mult_part_out08[410] <= P_11_8[31];
            mult_part_out08[411] <= P_15_6[12];
            mult_part_out08[412] <= P_12_7[40];
            mult_part_out08[413] <= P_14_6[31];
            mult_part_out08[414] <= P_13_8[1];
            mult_part_out08[415] <= P_10_9[29];
            mult_part_out08[416] <= P_11_8[37];
            mult_part_out08[417] <= P_13_8[4];
            mult_part_out08[418] <= P_11_9[15];
            mult_part_out08[419] <= P_13_8[6];
            mult_part_out08[420] <= P_14_7[14];
            mult_part_out08[421] <= P_10_9[35];
            mult_part_out08[422] <= P_10_9[36];
            mult_part_out08[423] <= P_15_6[24];
            mult_part_out08[424] <= P_13_7[35];
            mult_part_out08[425] <= P_12_9[5];
            mult_part_out08[426] <= P_14_7[20];
            mult_part_out08[427] <= P_10_10[17];
            mult_part_out08[428] <= P_12_8[32];
            mult_part_out08[429] <= P_13_7[40];
            mult_part_out08[430] <= P_12_9[10];
            mult_part_out08[431] <= P_14_7[25];
            mult_part_out08[432] <= P_14_7[26];
            mult_part_out08[433] <= P_11_9[30];
            mult_part_out08[434] <= P_10_10[24];
            mult_part_out08[435] <= P_11_10[8];
            mult_part_out08[436] <= P_14_8[6];
            mult_part_out08[437] <= P_11_10[10];
            mult_part_out08[438] <= P_10_10[28];
            mult_part_out08[439] <= P_13_9[2];
            mult_part_out08[440] <= P_10_10[30];
            mult_part_out08[441] <= P_10_10[31];
            mult_part_out08[442] <= P_14_7[36];

            mult_part_out09[96] <= P_0_3[24];
            mult_part_out09[97] <= P_0_3[25];
            mult_part_out09[98] <= P_0_4[2];
            mult_part_out09[99] <= P_0_4[3];
            mult_part_out09[100] <= P_0_3[28];
            mult_part_out09[101] <= P_3_1[26];
            mult_part_out09[102] <= P_0_3[30];
            mult_part_out09[103] <= P_0_4[7];
            mult_part_out09[104] <= P_3_2[5];
            mult_part_out09[105] <= P_3_1[30];
            mult_part_out09[106] <= P_0_3[34];
            mult_part_out09[107] <= P_3_2[8];
            mult_part_out09[108] <= P_2_2[26];
            mult_part_out09[109] <= P_3_2[10];
            mult_part_out09[110] <= P_5_1[1];
            mult_part_out09[111] <= P_5_1[2];
            mult_part_out09[112] <= P_5_1[3];
            mult_part_out09[113] <= P_1_4[0];
            mult_part_out09[114] <= P_1_3[25];
            mult_part_out09[115] <= P_5_0[30];
            mult_part_out09[116] <= P_2_2[34];
            mult_part_out09[117] <= P_6_0[15];
            mult_part_out09[118] <= P_6_0[16];
            mult_part_out09[119] <= P_4_1[27];
            mult_part_out09[120] <= P_3_2[21];
            mult_part_out09[121] <= P_6_0[19];
            mult_part_out09[122] <= P_2_3[16];
            mult_part_out09[123] <= P_0_5[3];
            mult_part_out09[124] <= P_3_3[1];
            mult_part_out09[125] <= P_1_3[36];
            mult_part_out09[126] <= P_1_3[37];
            mult_part_out09[127] <= P_6_1[1];
            mult_part_out09[128] <= P_6_0[26];
            mult_part_out09[129] <= P_1_3[40];
            mult_part_out09[130] <= P_4_2[14];
            mult_part_out09[131] <= P_6_1[5];
            mult_part_out09[132] <= P_6_0[30];
            mult_part_out09[133] <= P_2_4[3];
            mult_part_out09[134] <= P_3_2[35];
            mult_part_out09[135] <= P_4_2[19];
            mult_part_out09[136] <= P_6_0[34];
            mult_part_out09[137] <= P_6_0[35];
            mult_part_out09[138] <= P_1_4[25];
            mult_part_out09[139] <= P_2_3[33];
            mult_part_out09[140] <= P_2_3[34];
            mult_part_out09[141] <= P_5_2[8];
            mult_part_out09[142] <= P_7_0[23];
            mult_part_out09[143] <= P_5_2[10];
            mult_part_out09[144] <= P_1_5[7];
            mult_part_out09[145] <= P_2_3[39];
            mult_part_out09[146] <= P_8_0[10];
            mult_part_out09[147] <= P_6_1[21];
            mult_part_out09[148] <= P_1_4[35];
            mult_part_out09[149] <= P_7_0[30];
            mult_part_out09[150] <= P_0_5[30];
            mult_part_out09[151] <= P_1_4[38];
            mult_part_out09[152] <= P_6_1[26];
            mult_part_out09[153] <= P_9_0[0];
            mult_part_out09[154] <= P_1_5[17];
            mult_part_out09[155] <= P_3_3[32];
            mult_part_out09[156] <= P_4_3[16];
            mult_part_out09[157] <= P_0_5[37];
            mult_part_out09[158] <= P_4_3[18];
            mult_part_out09[159] <= P_0_5[39];
            mult_part_out09[160] <= P_4_3[20];
            mult_part_out09[161] <= P_6_2[11];
            mult_part_out09[162] <= P_5_2[29];
            mult_part_out09[163] <= P_6_2[13];
            mult_part_out09[164] <= P_4_3[24];
            mult_part_out09[165] <= P_2_5[11];
            mult_part_out09[166] <= P_6_1[40];
            mult_part_out09[167] <= P_8_1[7];
            mult_part_out09[168] <= P_7_1[25];
            mult_part_out09[169] <= P_4_4[5];
            mult_part_out09[170] <= P_0_6[26];
            mult_part_out09[171] <= P_7_2[4];
            mult_part_out09[172] <= P_8_1[12];
            mult_part_out09[173] <= P_6_2[23];
            mult_part_out09[174] <= P_5_3[17];
            mult_part_out09[175] <= P_6_2[25];
            mult_part_out09[176] <= P_1_5[39];
            mult_part_out09[177] <= P_2_5[23];
            mult_part_out09[178] <= P_7_2[11];
            mult_part_out09[179] <= P_4_3[39];
            mult_part_out09[180] <= P_0_7[12];
            mult_part_out09[181] <= P_7_2[14];
            mult_part_out09[182] <= P_8_1[22];
            mult_part_out09[183] <= P_7_2[16];
            mult_part_out09[184] <= P_5_3[27];
            mult_part_out09[185] <= P_9_1[8];
            mult_part_out09[186] <= P_6_2[36];
            mult_part_out09[187] <= P_6_2[37];
            mult_part_out09[188] <= P_1_6[27];
            mult_part_out09[189] <= P_9_0[36];
            mult_part_out09[190] <= P_1_7[5];
            mult_part_out09[191] <= P_3_5[20];
            mult_part_out09[192] <= P_7_3[1];
            mult_part_out09[193] <= P_7_3[2];
            mult_part_out09[194] <= P_7_3[3];
            mult_part_out09[195] <= P_10_0[25];
            mult_part_out09[196] <= P_1_7[11];
            mult_part_out09[197] <= P_1_7[12];
            mult_part_out09[198] <= P_3_6[3];
            mult_part_out09[199] <= P_11_0[12];
            mult_part_out09[200] <= P_5_4[19];
            mult_part_out09[201] <= P_1_7[16];
            mult_part_out09[202] <= P_2_6[24];
            mult_part_out09[203] <= P_3_5[32];
            mult_part_out09[204] <= P_0_8[12];
            mult_part_out09[205] <= P_12_0[1];
            mult_part_out09[206] <= P_9_1[29];
            mult_part_out09[207] <= P_1_7[22];
            mult_part_out09[208] <= P_12_0[4];
            mult_part_out09[209] <= P_1_7[24];
            mult_part_out09[210] <= P_1_7[25];
            mult_part_out09[211] <= P_5_4[30];
            mult_part_out09[212] <= P_9_2[11];
            mult_part_out09[213] <= P_11_1[2];
            mult_part_out09[214] <= P_8_2[30];
            mult_part_out09[215] <= P_5_4[34];
            mult_part_out09[216] <= P_10_1[22];
            mult_part_out09[217] <= P_7_3[26];
            mult_part_out09[218] <= P_7_3[27];
            mult_part_out09[219] <= P_0_8[27];
            mult_part_out09[220] <= P_8_2[36];
            mult_part_out09[221] <= P_0_9[5];
            mult_part_out09[222] <= P_10_1[28];
            mult_part_out09[223] <= P_1_8[14];
            mult_part_out09[224] <= P_4_5[36];
            mult_part_out09[225] <= P_11_0[38];
            mult_part_out09[226] <= P_6_5[4];
            mult_part_out09[227] <= P_1_8[18];
            mult_part_out09[228] <= P_2_7[26];
            mult_part_out09[229] <= P_6_4[31];
            mult_part_out09[230] <= P_9_3[5];
            mult_part_out09[231] <= P_12_0[27];
            mult_part_out09[232] <= P_11_1[21];
            mult_part_out09[233] <= P_9_3[8];
            mult_part_out09[234] <= P_3_7[15];
            mult_part_out09[235] <= P_3_6[40];
            mult_part_out09[236] <= P_3_7[17];
            mult_part_out09[237] <= P_13_0[16];
            mult_part_out09[238] <= P_7_4[23];
            mult_part_out09[239] <= P_1_8[30];
            mult_part_out09[240] <= P_7_4[25];
            mult_part_out09[241] <= P_8_4[9];
            mult_part_out09[242] <= P_10_2[24];
            mult_part_out09[243] <= P_2_8[17];
            mult_part_out09[244] <= P_14_0[6];
            mult_part_out09[245] <= P_3_8[2];
            mult_part_out09[246] <= P_12_1[18];
            mult_part_out09[247] <= P_6_5[25];
            mult_part_out09[248] <= P_4_7[12];
            mult_part_out09[249] <= P_12_1[21];
            mult_part_out09[250] <= P_4_7[14];
            mult_part_out09[251] <= P_3_7[32];
            mult_part_out09[252] <= P_4_7[16];
            mult_part_out09[253] <= P_13_1[8];
            mult_part_out09[254] <= P_9_3[29];
            mult_part_out09[255] <= P_5_6[26];
            mult_part_out09[256] <= P_12_1[28];
            mult_part_out09[257] <= P_10_3[15];
            mult_part_out09[258] <= P_3_8[15];
            mult_part_out09[259] <= P_2_8[33];
            mult_part_out09[260] <= P_13_1[15];
            mult_part_out09[261] <= P_14_0[23];
            mult_part_out09[262] <= P_2_8[36];
            mult_part_out09[263] <= P_12_1[35];
            mult_part_out09[264] <= P_2_8[38];
            mult_part_out09[265] <= P_2_9[15];
            mult_part_out09[266] <= P_1_9[33];
            mult_part_out09[267] <= P_8_4[35];
            mult_part_out09[268] <= P_4_7[32];
            mult_part_out09[269] <= P_6_6[23];
            mult_part_out09[270] <= P_5_7[17];
            mult_part_out09[271] <= P_12_2[19];
            mult_part_out09[272] <= P_15_0[17];
            mult_part_out09[273] <= P_12_2[21];
            mult_part_out09[274] <= P_11_3[15];
            mult_part_out09[275] <= P_10_3[33];
            mult_part_out09[276] <= P_2_10[2];
            mult_part_out09[277] <= P_10_4[11];
            mult_part_out09[278] <= P_6_7[8];
            mult_part_out09[279] <= P_2_10[5];
            mult_part_out09[280] <= P_14_1[18];
            mult_part_out09[281] <= P_2_10[7];
            mult_part_out09[282] <= P_4_8[22];
            mult_part_out09[283] <= P_5_8[6];
            mult_part_out09[284] <= P_13_2[15];
            mult_part_out09[285] <= P_11_3[26];
            mult_part_out09[286] <= P_14_1[24];
            mult_part_out09[287] <= P_14_1[25];
            mult_part_out09[288] <= P_4_9[4];
            mult_part_out09[289] <= P_1_10[32];
            mult_part_out09[290] <= P_11_4[7];
            mult_part_out09[291] <= P_10_4[25];
            mult_part_out09[292] <= P_15_1[13];
            mult_part_out09[293] <= P_7_6[30];
            mult_part_out09[294] <= P_3_10[3];
            mult_part_out09[295] <= P_2_10[21];
            mult_part_out09[296] <= P_11_3[37];
            mult_part_out09[297] <= P_13_3[4];
            mult_part_out09[298] <= P_7_6[35];
            mult_part_out09[299] <= P_8_6[19];
            mult_part_out09[300] <= P_12_3[24];
            mult_part_out09[301] <= P_12_3[25];
            mult_part_out09[302] <= P_6_8[8];
            mult_part_out09[303] <= P_9_6[6];
            mult_part_out09[304] <= P_14_2[18];
            mult_part_out09[305] <= P_3_10[14];
            mult_part_out09[306] <= P_10_4[40];
            mult_part_out09[307] <= P_8_6[27];
            mult_part_out09[308] <= P_8_7[4];
            mult_part_out09[309] <= P_13_3[16];
            mult_part_out09[310] <= P_4_9[26];
            mult_part_out09[311] <= P_14_2[25];
            mult_part_out09[312] <= P_15_2[9];
            mult_part_out09[313] <= P_15_2[10];
            mult_part_out09[314] <= P_8_6[34];
            mult_part_out09[315] <= P_14_2[29];
            mult_part_out09[316] <= P_6_8[22];
            mult_part_out09[317] <= P_4_10[9];
            mult_part_out09[318] <= P_5_9[17];
            mult_part_out09[319] <= P_6_8[25];
            mult_part_out09[320] <= P_8_7[16];
            mult_part_out09[321] <= P_7_8[10];
            mult_part_out09[322] <= P_13_3[29];
            mult_part_out09[323] <= P_6_8[29];
            mult_part_out09[324] <= P_9_6[27];
            mult_part_out09[325] <= P_7_7[38];
            mult_part_out09[326] <= P_7_7[39];
            mult_part_out09[327] <= P_11_5[20];
            mult_part_out09[328] <= P_12_5[4];
            mult_part_out09[329] <= P_9_6[32];
            mult_part_out09[330] <= P_11_5[23];
            mult_part_out09[331] <= P_9_6[34];
            mult_part_out09[332] <= P_13_4[15];
            mult_part_out09[333] <= P_9_7[12];
            mult_part_out09[334] <= P_11_6[3];
            mult_part_out09[335] <= P_4_10[27];
            mult_part_out09[336] <= P_11_6[5];
            mult_part_out09[337] <= P_5_10[12];
            mult_part_out09[338] <= P_15_3[11];
            mult_part_out09[339] <= P_7_8[28];
            mult_part_out09[340] <= P_8_8[12];
            mult_part_out09[341] <= P_10_7[3];
            mult_part_out09[342] <= P_13_4[25];
            mult_part_out09[343] <= P_8_7[39];
            mult_part_out09[344] <= P_12_5[20];
            mult_part_out09[345] <= P_13_5[4];
            mult_part_out09[346] <= P_14_3[36];
            mult_part_out09[347] <= P_9_7[26];
            mult_part_out09[348] <= P_11_6[17];
            mult_part_out09[349] <= P_12_6[1];
            mult_part_out09[350] <= P_6_10[8];
            mult_part_out09[351] <= P_10_6[37];
            mult_part_out09[352] <= P_6_10[10];
            mult_part_out09[353] <= P_12_6[5];
            mult_part_out09[354] <= P_8_8[26];
            mult_part_out09[355] <= P_12_6[7];
            mult_part_out09[356] <= P_6_9[38];
            mult_part_out09[357] <= P_8_9[5];
            mult_part_out09[358] <= P_13_5[17];
            mult_part_out09[359] <= P_10_7[21];
            mult_part_out09[360] <= P_15_4[9];
            mult_part_out09[361] <= P_14_5[3];
            mult_part_out09[362] <= P_11_6[31];
            mult_part_out09[363] <= P_6_10[21];
            mult_part_out09[364] <= P_13_5[23];
            mult_part_out09[365] <= P_6_10[23];
            mult_part_out09[366] <= P_8_9[14];
            mult_part_out09[367] <= P_15_4[16];
            mult_part_out09[368] <= P_12_6[20];
            mult_part_out09[369] <= P_11_6[38];
            mult_part_out09[370] <= P_9_8[25];
            mult_part_out09[371] <= P_7_9[36];
            mult_part_out09[372] <= P_10_8[10];
            mult_part_out09[373] <= P_9_9[4];
            mult_part_out09[374] <= P_13_5[33];
            mult_part_out09[375] <= P_9_8[30];
            mult_part_out09[376] <= P_10_7[38];
            mult_part_out09[377] <= P_14_5[19];
            mult_part_out09[378] <= P_13_6[13];
            mult_part_out09[379] <= P_7_10[20];
            mult_part_out09[380] <= P_9_8[35];
            mult_part_out09[381] <= P_12_7[9];
            mult_part_out09[382] <= P_8_10[6];
            mult_part_out09[383] <= P_8_10[7];
            mult_part_out09[384] <= P_9_9[15];
            mult_part_out09[385] <= P_9_8[40];
            mult_part_out09[386] <= P_12_6[38];
            mult_part_out09[387] <= P_15_5[12];
            mult_part_out09[388] <= P_9_9[19];
            mult_part_out09[389] <= P_13_6[24];
            mult_part_out09[390] <= P_7_10[31];
            mult_part_out09[391] <= P_11_7[36];
            mult_part_out09[392] <= P_10_8[30];
            mult_part_out09[393] <= P_9_9[24];
            mult_part_out09[394] <= P_10_9[8];
            mult_part_out09[395] <= P_13_6[30];
            mult_part_out09[396] <= P_13_7[7];
            mult_part_out09[397] <= P_9_9[28];
            mult_part_out09[398] <= P_9_10[5];
            mult_part_out09[399] <= P_14_6[17];
            mult_part_out09[400] <= P_9_9[31];
            mult_part_out09[401] <= P_13_7[12];
            mult_part_out09[402] <= P_13_7[13];
            mult_part_out09[403] <= P_9_10[10];
            mult_part_out09[404] <= P_12_8[8];
            mult_part_out09[405] <= P_15_6[6];
            mult_part_out09[406] <= P_11_8[27];
            mult_part_out09[407] <= P_12_8[11];
            mult_part_out09[408] <= P_14_6[26];
            mult_part_out09[409] <= P_10_9[23];
            mult_part_out09[410] <= P_9_10[17];
            mult_part_out09[411] <= P_12_7[39];
            mult_part_out09[412] <= P_13_7[23];
            mult_part_out09[413] <= P_15_6[14];
            mult_part_out09[414] <= P_10_9[28];
            mult_part_out09[415] <= P_14_7[9];
            mult_part_out09[416] <= P_13_8[3];
            mult_part_out09[417] <= P_10_10[7];
            mult_part_out09[418] <= P_9_10[25];
            mult_part_out09[419] <= P_14_7[13];
            mult_part_out09[420] <= P_13_8[7];
            mult_part_out09[421] <= P_13_7[32];
            mult_part_out09[422] <= P_15_6[23];
            mult_part_out09[423] <= P_15_7[0];
            mult_part_out09[424] <= P_10_9[38];
            mult_part_out09[425] <= P_15_7[2];

            mult_part_out10[102] <= P_4_1[10];
            mult_part_out10[103] <= P_5_0[18];
            mult_part_out10[104] <= P_1_2[39];
            mult_part_out10[105] <= P_4_1[13];
            mult_part_out10[106] <= P_4_1[14];
            mult_part_out10[107] <= P_5_0[22];
            mult_part_out10[108] <= P_3_2[9];
            mult_part_out10[109] <= P_6_0[7];
            mult_part_out10[110] <= P_0_4[14];
            mult_part_out10[111] <= P_2_3[5];
            mult_part_out10[112] <= P_2_3[6];
            mult_part_out10[113] <= P_3_2[14];
            mult_part_out10[114] <= P_3_2[15];
            mult_part_out10[115] <= P_3_2[16];
            mult_part_out10[116] <= P_2_3[10];
            mult_part_out10[117] <= P_3_2[18];
            mult_part_out10[118] <= P_2_2[36];
            mult_part_out10[119] <= P_3_2[20];
            mult_part_out10[120] <= P_6_0[18];
            mult_part_out10[121] <= P_0_5[1];
            mult_part_out10[122] <= P_4_2[6];
            mult_part_out10[123] <= P_1_3[34];
            mult_part_out10[124] <= P_4_1[32];
            mult_part_out10[125] <= P_0_4[29];
            mult_part_out10[126] <= P_3_3[3];
            mult_part_out10[127] <= P_4_2[11];
            mult_part_out10[128] <= P_1_4[15];
            mult_part_out10[129] <= P_4_2[13];
            mult_part_out10[130] <= P_5_1[21];
            mult_part_out10[131] <= P_4_2[15];
            mult_part_out10[132] <= P_0_5[12];
            mult_part_out10[133] <= P_7_0[14];
            mult_part_out10[134] <= P_0_5[14];
            mult_part_out10[135] <= P_2_4[5];
            mult_part_out10[136] <= P_0_4[40];
            mult_part_out10[137] <= P_2_4[7];
            mult_part_out10[138] <= P_3_2[39];
            mult_part_out10[139] <= P_4_2[23];
            mult_part_out10[140] <= P_5_1[31];
            mult_part_out10[141] <= P_6_1[15];
            mult_part_out10[142] <= P_5_1[33];
            mult_part_out10[143] <= P_2_3[37];
            mult_part_out10[144] <= P_5_2[11];
            mult_part_out10[145] <= P_7_1[2];
            mult_part_out10[146] <= P_4_3[6];
            mult_part_out10[147] <= P_0_6[3];
            mult_part_out10[148] <= P_4_3[8];
            mult_part_out10[149] <= P_8_0[13];
            mult_part_out10[150] <= P_4_3[10];
            mult_part_out10[151] <= P_7_1[8];
            mult_part_out10[152] <= P_2_4[22];
            mult_part_out10[153] <= P_7_1[10];
            mult_part_out10[154] <= P_4_3[14];
            mult_part_out10[155] <= P_2_5[1];
            mult_part_out10[156] <= P_6_2[6];
            mult_part_out10[157] <= P_1_5[20];
            mult_part_out10[158] <= P_7_1[15];
            mult_part_out10[159] <= P_6_1[33];
            mult_part_out10[160] <= P_8_1[0];
            mult_part_out10[161] <= P_3_3[38];
            mult_part_out10[162] <= P_3_3[39];
            mult_part_out10[163] <= P_6_1[37];
            mult_part_out10[164] <= P_6_1[38];
            mult_part_out10[165] <= P_8_0[29];
            mult_part_out10[166] <= P_3_4[19];
            mult_part_out10[167] <= P_2_5[13];
            mult_part_out10[168] <= P_5_2[35];
            mult_part_out10[169] <= P_1_5[32];
            mult_part_out10[170] <= P_1_5[33];
            mult_part_out10[171] <= P_7_1[28];
            mult_part_out10[172] <= P_8_0[36];
            mult_part_out10[173] <= P_0_7[5];
            mult_part_out10[174] <= P_6_2[24];
            mult_part_out10[175] <= P_4_3[35];
            mult_part_out10[176] <= P_5_3[19];
            mult_part_out10[177] <= P_6_2[27];
            mult_part_out10[178] <= P_10_0[8];
            mult_part_out10[179] <= P_9_1[2];
            mult_part_out10[180] <= P_9_1[3];
            mult_part_out10[181] <= P_4_4[17];
            mult_part_out10[182] <= P_9_1[5];
            mult_part_out10[183] <= P_4_4[19];
            mult_part_out10[184] <= P_9_1[7];
            mult_part_out10[185] <= P_7_2[18];
            mult_part_out10[186] <= P_2_6[8];
            mult_part_out10[187] <= P_8_2[3];
            mult_part_out10[188] <= P_2_5[34];
            mult_part_out10[189] <= P_6_2[39];
            mult_part_out10[190] <= P_9_1[13];
            mult_part_out10[191] <= P_9_0[38];
            mult_part_out10[192] <= P_3_5[21];
            mult_part_out10[193] <= P_6_3[19];
            mult_part_out10[194] <= P_1_6[33];
            mult_part_out10[195] <= P_5_3[38];
            mult_part_out10[196] <= P_3_6[1];
            mult_part_out10[197] <= P_4_5[9];
            mult_part_out10[198] <= P_5_4[17];
            mult_part_out10[199] <= P_7_3[8];
            mult_part_out10[200] <= P_0_7[32];
            mult_part_out10[201] <= P_2_6[23];
            mult_part_out10[202] <= P_0_7[34];
            mult_part_out10[203] <= P_2_7[1];
            mult_part_out10[204] <= P_3_5[33];
            mult_part_out10[205] <= P_7_2[38];
            mult_part_out10[206] <= P_4_5[18];
            mult_part_out10[207] <= P_3_5[36];
            mult_part_out10[208] <= P_5_4[27];
            mult_part_out10[209] <= P_11_0[22];
            mult_part_out10[210] <= P_2_6[32];
            mult_part_out10[211] <= P_6_4[13];
            mult_part_out10[212] <= P_4_5[24];
            mult_part_out10[213] <= P_6_4[15];
            mult_part_out10[214] <= P_3_6[19];
            mult_part_out10[215] <= P_8_3[7];
            mult_part_out10[216] <= P_7_3[25];
            mult_part_out10[217] <= P_2_7[15];
            mult_part_out10[218] <= P_11_0[31];
            mult_part_out10[219] <= P_4_5[31];
            mult_part_out10[220] <= P_3_6[25];
            mult_part_out10[221] <= P_11_0[34];
            mult_part_out10[222] <= P_11_1[11];
            mult_part_out10[223] <= P_6_5[1];
            mult_part_out10[224] <= P_7_3[33];
            mult_part_out10[225] <= P_9_2[24];
            mult_part_out10[226] <= P_9_2[25];
            mult_part_out10[227] <= P_5_5[22];
            mult_part_out10[228] <= P_7_3[37];
            mult_part_out10[229] <= P_13_0[8];
            mult_part_out10[230] <= P_9_2[29];
            mult_part_out10[231] <= P_7_3[40];
            mult_part_out10[232] <= P_12_0[28];
            mult_part_out10[233] <= P_3_7[14];
            mult_part_out10[234] <= P_3_6[39];
            mult_part_out10[235] <= P_2_8[9];
            mult_part_out10[236] <= P_6_5[14];
            mult_part_out10[237] <= P_12_0[33];
            mult_part_out10[238] <= P_12_1[10];
            mult_part_out10[239] <= P_14_0[1];
            mult_part_out10[240] <= P_8_4[8];
            mult_part_out10[241] <= P_7_5[2];
            mult_part_out10[242] <= P_0_10[2];
            mult_part_out10[243] <= P_3_8[0];
            mult_part_out10[244] <= P_4_7[8];
            mult_part_out10[245] <= P_8_3[37];
            mult_part_out10[246] <= P_13_0[25];
            mult_part_out10[247] <= P_0_9[31];
            mult_part_out10[248] <= P_13_0[27];
            mult_part_out10[249] <= P_9_3[24];
            mult_part_out10[250] <= P_6_6[4];
            mult_part_out10[251] <= P_11_2[16];
            mult_part_out10[252] <= P_10_2[34];
            mult_part_out10[253] <= P_12_1[25];
            mult_part_out10[254] <= P_7_5[15];
            mult_part_out10[255] <= P_13_1[10];
            mult_part_out10[256] <= P_6_5[34];
            mult_part_out10[257] <= P_8_5[1];
            mult_part_out10[258] <= P_9_4[9];
            mult_part_out10[259] <= P_0_10[19];
            mult_part_out10[260] <= P_14_0[22];
            mult_part_out10[261] <= P_3_8[18];
            mult_part_out10[262] <= P_13_1[17];
            mult_part_out10[263] <= P_14_0[25];
            mult_part_out10[264] <= P_12_1[36];
            mult_part_out10[265] <= P_9_3[40];
            mult_part_out10[266] <= P_1_10[9];
            mult_part_out10[267] <= P_13_1[22];
            mult_part_out10[268] <= P_11_3[9];
            mult_part_out10[269] <= P_3_8[26];
            mult_part_out10[270] <= P_1_10[13];
            mult_part_out10[271] <= P_13_1[26];
            mult_part_out10[272] <= P_2_9[22];
            mult_part_out10[273] <= P_14_1[11];
            mult_part_out10[274] <= P_4_7[38];
            mult_part_out10[275] <= P_9_5[2];
            mult_part_out10[276] <= P_6_6[30];
            mult_part_out10[277] <= P_2_9[27];
            mult_part_out10[278] <= P_14_0[40];
            mult_part_out10[279] <= P_7_6[16];
            mult_part_out10[280] <= P_3_9[13];
            mult_part_out10[281] <= P_10_4[15];
            mult_part_out10[282] <= P_9_5[9];
            mult_part_out10[283] <= P_11_4[0];
            mult_part_out10[284] <= P_2_10[10];
            mult_part_out10[285] <= P_14_1[23];
            mult_part_out10[286] <= P_8_6[6];
            mult_part_out10[287] <= P_9_5[14];
            mult_part_out10[288] <= P_15_1[9];
            mult_part_out10[289] <= P_3_9[22];
            mult_part_out10[290] <= P_4_9[6];
            mult_part_out10[291] <= P_7_6[28];
            mult_part_out10[292] <= P_4_8[32];
            mult_part_out10[293] <= P_14_2[7];
            mult_part_out10[294] <= P_6_8[0];
            mult_part_out10[295] <= P_4_8[35];
            mult_part_out10[296] <= P_13_2[27];
            mult_part_out10[297] <= P_8_6[17];
            mult_part_out10[298] <= P_11_4[15];
            mult_part_out10[299] <= P_12_3[23];
            mult_part_out10[300] <= P_5_8[23];
            mult_part_out10[301] <= P_14_2[15];
            mult_part_out10[302] <= P_7_7[15];
            mult_part_out10[303] <= P_15_1[24];
            mult_part_out10[304] <= P_3_9[37];
            mult_part_out10[305] <= P_5_9[4];
            mult_part_out10[306] <= P_14_2[20];
            mult_part_out10[307] <= P_6_7[37];
            mult_part_out10[308] <= P_11_4[25];
            mult_part_out10[309] <= P_11_5[2];
            mult_part_out10[310] <= P_10_5[20];
            mult_part_out10[311] <= P_4_10[3];
            mult_part_out10[312] <= P_5_9[11];
            mult_part_out10[313] <= P_13_3[20];
            mult_part_out10[314] <= P_5_9[13];
            mult_part_out10[315] <= P_7_7[28];
            mult_part_out10[316] <= P_9_6[19];
            mult_part_out10[317] <= P_3_10[26];
            mult_part_out10[318] <= P_12_4[18];
            mult_part_out10[319] <= P_7_8[8];
            mult_part_out10[320] <= P_6_9[2];
            mult_part_out10[321] <= P_4_9[37];
            mult_part_out10[322] <= P_10_5[32];
            mult_part_out10[323] <= P_9_7[2];
            mult_part_out10[324] <= P_7_7[37];
            mult_part_out10[325] <= P_4_10[17];
            mult_part_out10[326] <= P_4_10[18];
            mult_part_out10[327] <= P_7_8[16];
            mult_part_out10[328] <= P_9_6[31];
            mult_part_out10[329] <= P_10_6[15];
            mult_part_out10[330] <= P_5_9[29];
            mult_part_out10[331] <= P_7_8[20];
            mult_part_out10[332] <= P_12_4[32];
            mult_part_out10[333] <= P_11_6[2];
            mult_part_out10[334] <= P_12_4[34];
            mult_part_out10[335] <= P_6_9[17];
            mult_part_out10[336] <= P_7_9[1];
            mult_part_out10[337] <= P_9_6[40];
            mult_part_out10[338] <= P_8_8[10];
            mult_part_out10[339] <= P_10_6[25];
            mult_part_out10[340] <= P_12_5[16];
            mult_part_out10[341] <= P_8_8[13];
            mult_part_out10[342] <= P_8_7[38];
            mult_part_out10[343] <= P_6_10[1];
            mult_part_out10[344] <= P_10_6[30];
            mult_part_out10[345] <= P_9_7[24];
            mult_part_out10[346] <= P_7_9[11];
            mult_part_out10[347] <= P_9_8[2];
            mult_part_out10[348] <= P_7_8[37];
            mult_part_out10[349] <= P_14_4[15];
            mult_part_out10[350] <= P_7_8[39];
            mult_part_out10[351] <= P_11_6[20];
            mult_part_out10[352] <= P_11_6[21];
            mult_part_out10[353] <= P_9_8[8];
            mult_part_out10[354] <= P_12_5[30];
            mult_part_out10[355] <= P_6_10[13];
            mult_part_out10[356] <= P_13_4[39];
            mult_part_out10[357] <= P_6_9[39];
            mult_part_out10[358] <= P_14_5[0];
            mult_part_out10[359] <= P_12_5[35];
            mult_part_out10[360] <= P_12_5[36];
            mult_part_out10[361] <= P_12_6[13];
            mult_part_out10[362] <= P_15_4[11];
            mult_part_out10[363] <= P_9_8[18];
            mult_part_out10[364] <= P_7_9[29];
            mult_part_out10[365] <= P_14_5[7];
            mult_part_out10[366] <= P_7_10[7];
            mult_part_out10[367] <= P_14_5[9];
            mult_part_out10[368] <= P_13_5[27];
            mult_part_out10[369] <= P_14_5[11];
            mult_part_out10[370] <= P_11_7[15];
            mult_part_out10[371] <= P_13_5[30];
            mult_part_out10[372] <= P_9_9[3];
            mult_part_out10[373] <= P_10_7[35];
            mult_part_out10[374] <= P_11_7[19];
            mult_part_out10[375] <= P_10_8[13];
            mult_part_out10[376] <= P_11_7[21];
            mult_part_out10[377] <= P_10_8[15];
            mult_part_out10[378] <= P_13_5[37];
            mult_part_out10[379] <= P_9_8[34];
            mult_part_out10[380] <= P_11_8[1];
            mult_part_out10[381] <= P_12_6[33];
            mult_part_out10[382] <= P_11_8[3];
            mult_part_out10[383] <= P_14_6[1];
            mult_part_out10[384] <= P_8_9[32];
            mult_part_out10[385] <= P_9_9[16];
            mult_part_out10[386] <= P_8_9[34];
            mult_part_out10[387] <= P_10_8[25];
            mult_part_out10[388] <= P_11_7[33];
            mult_part_out10[389] <= P_14_6[7];
            mult_part_out10[390] <= P_9_9[21];
            mult_part_out10[391] <= P_14_6[9];
            mult_part_out10[392] <= P_13_7[3];
            mult_part_out10[393] <= P_11_7[38];
            mult_part_out10[394] <= P_9_10[1];
            mult_part_out10[395] <= P_10_8[33];
            mult_part_out10[396] <= P_14_6[14];
            mult_part_out10[397] <= P_9_10[4];
            mult_part_out10[398] <= P_10_8[36];
            mult_part_out10[399] <= P_13_6[34];
            mult_part_out10[400] <= P_12_7[28];
            mult_part_out10[401] <= P_12_8[5];
            mult_part_out10[402] <= P_9_9[33];
            mult_part_out10[403] <= P_13_7[14];
            mult_part_out10[404] <= P_13_7[15];
            mult_part_out10[405] <= P_11_8[26];
            mult_part_out10[406] <= P_8_10[30];
            mult_part_out10[407] <= P_13_7[18];
            mult_part_out10[408] <= P_9_10[15];
            mult_part_out10[409] <= P_11_8[30];
            mult_part_out10[410] <= P_14_6[28];
            mult_part_out10[411] <= P_10_10[1];
            mult_part_out10[412] <= P_10_9[26];
            mult_part_out10[413] <= P_10_9[27];
            mult_part_out10[414] <= P_14_7[8];
            mult_part_out10[415] <= P_9_10[22];
            mult_part_out10[416] <= P_15_6[17];
            mult_part_out10[417] <= P_11_8[38];
            mult_part_out10[418] <= P_14_6[36];
            mult_part_out10[419] <= P_11_9[16];
            mult_part_out10[420] <= P_10_9[34];
            mult_part_out10[421] <= P_10_10[11];
            mult_part_out10[422] <= P_9_10[29];
            mult_part_out10[423] <= P_13_8[10];

            mult_part_out11[119] <= P_7_0[0];
            mult_part_out11[120] <= P_0_5[0];
            mult_part_out11[121] <= P_5_1[12];
            mult_part_out11[122] <= P_2_2[40];
            mult_part_out11[123] <= P_3_3[0];
            mult_part_out11[124] <= P_5_1[15];
            mult_part_out11[125] <= P_5_1[16];
            mult_part_out11[126] <= P_6_0[24];
            mult_part_out11[127] <= P_1_3[38];
            mult_part_out11[128] <= P_4_2[12];
            mult_part_out11[129] <= P_3_3[6];
            mult_part_out11[130] <= P_3_3[7];
            mult_part_out11[131] <= P_4_1[39];
            mult_part_out11[132] <= P_3_2[33];
            mult_part_out11[133] <= P_4_2[17];
            mult_part_out11[134] <= P_5_1[25];
            mult_part_out11[135] <= P_6_1[9];
            mult_part_out11[136] <= P_2_3[30];
            mult_part_out11[137] <= P_4_2[21];
            mult_part_out11[138] <= P_8_0[2];
            mult_part_out11[139] <= P_3_2[40];
            mult_part_out11[140] <= P_7_0[21];
            mult_part_out11[141] <= P_0_5[21];
            mult_part_out11[142] <= P_1_5[5];
            mult_part_out11[143] <= P_8_0[7];
            mult_part_out11[144] <= P_7_1[1];
            mult_part_out11[145] <= P_5_2[12];
            mult_part_out11[146] <= P_0_6[2];
            mult_part_out11[147] <= P_4_3[7];
            mult_part_out11[148] <= P_2_4[18];
            mult_part_out11[149] <= P_1_4[36];
            mult_part_out11[150] <= P_1_5[13];
            mult_part_out11[151] <= P_6_1[25];
            mult_part_out11[152] <= P_4_2[36];
            mult_part_out11[153] <= P_3_3[30];
            mult_part_out11[154] <= P_9_0[1];
            mult_part_out11[155] <= P_0_5[35];
            mult_part_out11[156] <= P_1_5[19];
            mult_part_out11[157] <= P_2_4[27];
            mult_part_out11[158] <= P_2_5[4];
            mult_part_out11[159] <= P_5_2[26];
            mult_part_out11[160] <= P_5_3[3];
            mult_part_out11[161] <= P_2_4[31];
            mult_part_out11[162] <= P_6_2[12];
            mult_part_out11[163] <= P_9_0[10];
            mult_part_out11[164] <= P_0_6[20];
            mult_part_out11[165] <= P_1_6[4];
            mult_part_out11[166] <= P_4_4[2];
            mult_part_out11[167] <= P_8_0[31];
            mult_part_out11[168] <= P_2_5[14];
            mult_part_out11[169] <= P_1_6[8];
            mult_part_out11[170] <= P_5_3[13];
            mult_part_out11[171] <= P_1_6[10];
            mult_part_out11[172] <= P_4_3[32];
            mult_part_out11[173] <= P_3_4[26];
            mult_part_out11[174] <= P_9_0[21];
            mult_part_out11[175] <= P_7_1[32];
            mult_part_out11[176] <= P_10_0[6];
            mult_part_out11[177] <= P_4_3[37];
            mult_part_out11[178] <= P_9_0[25];
            mult_part_out11[179] <= P_9_0[26];
            mult_part_out11[180] <= P_5_3[23];
            mult_part_out11[181] <= P_5_4[0];
            mult_part_out11[182] <= P_6_2[32];
            mult_part_out11[183] <= P_10_0[13];
            mult_part_out11[184] <= P_9_0[31];
            mult_part_out11[185] <= P_6_3[11];
            mult_part_out11[186] <= P_4_4[22];
            mult_part_out11[187] <= P_2_6[9];
            mult_part_out11[188] <= P_1_7[3];
            mult_part_out11[189] <= P_0_7[21];
            mult_part_out11[190] <= P_2_6[12];
            mult_part_out11[191] <= P_1_6[30];
            mult_part_out11[192] <= P_6_3[18];
            mult_part_out11[193] <= P_5_4[12];
            mult_part_out11[194] <= P_0_7[26];
            mult_part_out11[195] <= P_3_5[24];
            mult_part_out11[196] <= P_3_5[25];
            mult_part_out11[197] <= P_0_7[29];
            mult_part_out11[198] <= P_3_5[27];
            mult_part_out11[199] <= P_6_3[25];
            mult_part_out11[200] <= P_8_1[40];
            mult_part_out11[201] <= P_3_5[30];
            mult_part_out11[202] <= P_11_0[15];
            mult_part_out11[203] <= P_2_6[25];
            mult_part_out11[204] <= P_10_0[34];
            mult_part_out11[205] <= P_5_5[0];
            mult_part_out11[206] <= P_2_6[28];
            mult_part_out11[207] <= P_4_5[19];
            mult_part_out11[208] <= P_1_7[23];
            mult_part_out11[209] <= P_9_1[32];
            mult_part_out11[210] <= P_3_5[39];
            mult_part_out11[211] <= P_2_6[33];
            mult_part_out11[212] <= P_2_6[34];
            mult_part_out11[213] <= P_10_1[19];
            mult_part_out11[214] <= P_12_0[10];
            mult_part_out11[215] <= P_9_1[38];
            mult_part_out11[216] <= P_9_2[15];
            mult_part_out11[217] <= P_12_0[13];
            mult_part_out11[218] <= P_2_6[40];
            mult_part_out11[219] <= P_10_2[1];
            mult_part_out11[220] <= P_10_1[26];
            mult_part_out11[221] <= P_1_7[36];
            mult_part_out11[222] <= P_7_4[7];
            mult_part_out11[223] <= P_10_2[5];
            mult_part_out11[224] <= P_9_2[23];
            mult_part_out11[225] <= P_4_5[37];
            mult_part_out11[226] <= P_7_4[11];
            mult_part_out11[227] <= P_10_1[33];
            mult_part_out11[228] <= P_9_3[3];
            mult_part_out11[229] <= P_3_6[34];
            mult_part_out11[230] <= P_7_3[39];
            mult_part_out11[231] <= P_7_4[16];
            mult_part_out11[232] <= P_9_3[7];
            mult_part_out11[233] <= P_12_0[29];
            mult_part_out11[234] <= P_12_0[30];
            mult_part_out11[235] <= P_1_9[2];
            mult_part_out11[236] <= P_4_7[0];
            mult_part_out11[237] <= P_8_3[29];
            mult_part_out11[238] <= P_4_7[2];
            mult_part_out11[239] <= P_0_9[23];
            mult_part_out11[240] <= P_3_7[21];
            mult_part_out11[241] <= P_0_10[1];
            mult_part_out11[242] <= P_2_8[16];
            mult_part_out11[243] <= P_5_5[38];
            mult_part_out11[244] <= P_10_3[2];
            mult_part_out11[245] <= P_6_5[23];
            mult_part_out11[246] <= P_1_8[37];
            mult_part_out11[247] <= P_3_7[28];
            mult_part_out11[248] <= P_1_8[39];
            mult_part_out11[249] <= P_0_10[9];
            mult_part_out11[250] <= P_12_1[22];
            mult_part_out11[251] <= P_4_7[15];
            mult_part_out11[252] <= P_6_5[30];
            mult_part_out11[253] <= P_2_8[27];
            mult_part_out11[254] <= P_0_9[38];
            mult_part_out11[255] <= P_12_1[27];
            mult_part_out11[256] <= P_9_4[7];
            mult_part_out11[257] <= P_5_6[28];
            mult_part_out11[258] <= P_10_3[16];
            mult_part_out11[259] <= P_6_5[37];
            mult_part_out11[260] <= P_9_3[35];
            mult_part_out11[261] <= P_1_10[4];
            mult_part_out11[262] <= P_2_9[12];
            mult_part_out11[263] <= P_15_0[8];
            mult_part_out11[264] <= P_4_8[4];
            mult_part_out11[265] <= P_10_3[23];
            mult_part_out11[266] <= P_8_5[10];
            mult_part_out11[267] <= P_7_6[4];
            mult_part_out11[268] <= P_5_7[15];
            mult_part_out11[269] <= P_2_9[19];
            mult_part_out11[270] <= P_4_8[10];
            mult_part_out11[271] <= P_4_7[35];
            mult_part_out11[272] <= P_4_7[36];
            mult_part_out11[273] <= P_6_7[3];
            mult_part_out11[274] <= P_13_2[5];
            mult_part_out11[275] <= P_14_1[13];
            mult_part_out11[276] <= P_14_0[38];
            mult_part_out11[277] <= P_12_2[25];
            mult_part_out11[278] <= P_5_7[25];
            mult_part_out11[279] <= P_5_8[2];
            mult_part_out11[280] <= P_1_10[23];
            mult_part_out11[281] <= P_9_4[32];
            mult_part_out11[282] <= P_5_7[29];
            mult_part_out11[283] <= P_12_2[31];
            mult_part_out11[284] <= P_14_1[22];
            mult_part_out11[285] <= P_12_3[9];
            mult_part_out11[286] <= P_9_5[13];
            mult_part_out11[287] <= P_13_2[18];
            mult_part_out11[288] <= P_1_10[31];
            mult_part_out11[289] <= P_6_7[19];
            mult_part_out11[290] <= P_5_7[37];
            mult_part_out11[291] <= P_11_4[8];
            mult_part_out11[292] <= P_5_7[39];
            mult_part_out11[293] <= P_5_7[40];
            mult_part_out11[294] <= P_10_5[4];
            mult_part_out11[295] <= P_6_7[25];
            mult_part_out11[296] <= P_4_8[36];
            mult_part_out11[297] <= P_7_7[10];
            mult_part_out11[298] <= P_9_6[1];
            mult_part_out11[299] <= P_9_5[26];
            mult_part_out11[300] <= P_4_9[16];
            mult_part_out11[301] <= P_7_6[38];
            mult_part_out11[302] <= P_2_10[28];
            mult_part_out11[303] <= P_3_10[12];
            mult_part_out11[304] <= P_5_8[27];
            mult_part_out11[305] <= P_8_7[1];
            mult_part_out11[306] <= P_3_9[39];
            mult_part_out11[307] <= P_3_10[16];
            mult_part_out11[308] <= P_9_5[35];
            mult_part_out11[309] <= P_13_2[40];
            mult_part_out11[310] <= P_5_9[9];
            mult_part_out11[311] <= P_11_4[28];
            mult_part_out11[312] <= P_8_6[32];
            mult_part_out11[313] <= P_5_8[36];
            mult_part_out11[314] <= P_12_3[38];
            mult_part_out11[315] <= P_12_3[39];
            mult_part_out11[316] <= P_14_3[6];
            mult_part_out11[317] <= P_5_9[16];
            mult_part_out11[318] <= P_6_8[24];
            mult_part_out11[319] <= P_8_6[39];
            mult_part_out11[320] <= P_10_6[6];
            mult_part_out11[321] <= P_15_2[18];
            mult_part_out11[322] <= P_5_9[21];
            mult_part_out11[323] <= P_4_9[39];
            mult_part_out11[324] <= P_4_10[16];
            mult_part_out11[325] <= P_13_3[32];
            mult_part_out11[326] <= P_13_3[33];
            mult_part_out11[327] <= P_13_3[34];
            mult_part_out11[328] <= P_9_7[7];
            mult_part_out11[329] <= P_14_3[19];
            mult_part_out11[330] <= P_12_5[6];
            mult_part_out11[331] <= P_4_10[23];
            mult_part_out11[332] <= P_7_8[21];
            mult_part_out11[333] <= P_12_5[9];
            mult_part_out11[334] <= P_6_9[16];
            mult_part_out11[335] <= P_9_7[14];
            mult_part_out11[336] <= P_4_10[28];
            mult_part_out11[337] <= P_11_5[30];
            mult_part_out11[338] <= P_4_10[30];
            mult_part_out11[339] <= P_10_7[1];
            mult_part_out11[340] <= P_4_10[32];
            mult_part_out11[341] <= P_10_6[27];
            mult_part_out11[342] <= P_14_3[32];
            mult_part_out11[343] <= P_7_9[8];
            mult_part_out11[344] <= P_7_8[33];
            mult_part_out11[345] <= P_9_8[0];
            mult_part_out11[346] <= P_10_6[32];
            mult_part_out11[347] <= P_14_3[37];
            mult_part_out11[348] <= P_15_3[21];
            mult_part_out11[349] <= P_13_5[8];
            mult_part_out11[350] <= P_12_5[26];
            mult_part_out11[351] <= P_6_9[33];
            mult_part_out11[352] <= P_6_9[34];
            mult_part_out11[353] <= P_11_6[22];
            mult_part_out11[354] <= P_12_6[6];
            mult_part_out11[355] <= P_14_4[21];
            mult_part_out11[356] <= P_8_9[4];
            mult_part_out11[357] <= P_5_10[32];
            mult_part_out11[358] <= P_12_5[34];
            mult_part_out11[359] <= P_8_9[7];
            mult_part_out11[360] <= P_11_6[29];
            mult_part_out11[361] <= P_7_10[2];
            mult_part_out11[362] <= P_9_8[17];
            mult_part_out11[363] <= P_7_9[28];
            mult_part_out11[364] <= P_10_8[2];
            mult_part_out11[365] <= P_10_7[27];
            mult_part_out11[366] <= P_11_7[11];
            mult_part_out11[367] <= P_10_7[29];
            mult_part_out11[368] <= P_13_6[3];
            mult_part_out11[369] <= P_14_4[35];
            mult_part_out11[370] <= P_8_9[18];
            mult_part_out11[371] <= P_6_10[29];
            mult_part_out11[372] <= P_7_10[13];
            mult_part_out11[373] <= P_11_7[18];
            mult_part_out11[374] <= P_9_8[29];
            mult_part_out11[375] <= P_15_4[24];
            mult_part_out11[376] <= P_9_9[7];
            mult_part_out11[377] <= P_12_7[5];
            mult_part_out11[378] <= P_12_6[30];
            mult_part_out11[379] <= P_9_9[10];
            mult_part_out11[380] <= P_13_6[15];
            mult_part_out11[381] <= P_8_9[29];
            mult_part_out11[382] <= P_8_9[30];
            mult_part_out11[383] <= P_12_7[11];
            mult_part_out11[384] <= P_14_6[2];
            mult_part_out11[385] <= P_12_7[13];
            mult_part_out11[386] <= P_14_5[28];
            mult_part_out11[387] <= P_13_6[22];
            mult_part_out11[388] <= P_8_9[36];
            mult_part_out11[389] <= P_10_8[27];
            mult_part_out11[390] <= P_10_8[28];
            mult_part_out11[391] <= P_13_6[26];
            mult_part_out11[392] <= P_9_9[23];
            mult_part_out11[393] <= P_13_7[4];
            mult_part_out11[394] <= P_13_7[5];
            mult_part_out11[395] <= P_14_6[13];
            mult_part_out11[396] <= P_10_9[10];
            mult_part_out11[397] <= P_12_8[1];
            mult_part_out11[398] <= P_8_10[22];
            mult_part_out11[399] <= P_12_7[27];
            mult_part_out11[400] <= P_15_6[1];
            mult_part_out11[401] <= P_8_10[25];
            mult_part_out11[402] <= P_12_7[30];
            mult_part_out11[403] <= P_10_9[17];
            mult_part_out11[404] <= P_11_9[1];
            mult_part_out11[405] <= P_11_9[2];
            mult_part_out11[406] <= P_12_7[34];
            mult_part_out11[407] <= P_14_6[25];
            mult_part_out11[408] <= P_14_7[2];

            mult_part_out12[120] <= P_4_2[4];
            mult_part_out12[121] <= P_3_2[22];
            mult_part_out12[122] <= P_1_3[33];
            mult_part_out12[123] <= P_7_0[4];
            mult_part_out12[124] <= P_3_2[25];
            mult_part_out12[125] <= P_3_3[2];
            mult_part_out12[126] <= P_4_1[34];
            mult_part_out12[127] <= P_3_3[4];
            mult_part_out12[128] <= P_3_3[5];
            mult_part_out12[129] <= P_1_4[16];
            mult_part_out12[130] <= P_1_4[17];
            mult_part_out12[131] <= P_3_3[8];
            mult_part_out12[132] <= P_4_1[40];
            mult_part_out12[133] <= P_0_4[37];
            mult_part_out12[134] <= P_6_0[32];
            mult_part_out12[135] <= P_6_0[33];
            mult_part_out12[136] <= P_2_4[6];
            mult_part_out12[137] <= P_2_3[31];
            mult_part_out12[138] <= P_4_2[22];
            mult_part_out12[139] <= P_0_5[19];
            mult_part_out12[140] <= P_6_0[38];
            mult_part_out12[141] <= P_3_3[18];
            mult_part_out12[142] <= P_1_4[29];
            mult_part_out12[143] <= P_6_1[17];
            mult_part_out12[144] <= P_4_2[28];
            mult_part_out12[145] <= P_6_1[19];
            mult_part_out12[146] <= P_7_1[3];
            mult_part_out12[147] <= P_5_2[14];
            mult_part_out12[148] <= P_0_6[4];
            mult_part_out12[149] <= P_7_1[6];
            mult_part_out12[150] <= P_0_6[6];
            mult_part_out12[151] <= P_5_2[18];
            mult_part_out12[152] <= P_3_3[29];
            mult_part_out12[153] <= P_6_1[27];
            mult_part_out12[154] <= P_3_3[31];
            mult_part_out12[155] <= P_1_5[18];
            mult_part_out12[156] <= P_7_1[13];
            mult_part_out12[157] <= P_5_2[24];
            mult_part_out12[158] <= P_9_0[5];
            mult_part_out12[159] <= P_0_6[15];
            mult_part_out12[160] <= P_2_4[30];
            mult_part_out12[161] <= P_8_1[1];
            mult_part_out12[162] <= P_8_1[2];
            mult_part_out12[163] <= P_0_6[19];
            mult_part_out12[164] <= P_2_4[34];
            mult_part_out12[165] <= P_6_2[15];
            mult_part_out12[166] <= P_9_0[13];
            mult_part_out12[167] <= P_7_1[24];
            mult_part_out12[168] <= P_0_6[24];
            mult_part_out12[169] <= P_6_2[19];
            mult_part_out12[170] <= P_8_0[34];
            mult_part_out12[171] <= P_3_5[0];
            mult_part_out12[172] <= P_5_2[39];
            mult_part_out12[173] <= P_5_3[16];
            mult_part_out12[174] <= P_10_0[4];
            mult_part_out12[175] <= P_3_4[28];
            mult_part_out12[176] <= P_3_5[5];
            mult_part_out12[177] <= P_0_6[33];
            mult_part_out12[178] <= P_4_3[38];
            mult_part_out12[179] <= P_8_1[19];
            mult_part_out12[180] <= P_4_4[16];
            mult_part_out12[181] <= P_2_6[3];
            mult_part_out12[182] <= P_7_1[39];
            mult_part_out12[183] <= P_5_4[2];
            mult_part_out12[184] <= P_2_6[6];
            mult_part_out12[185] <= P_4_4[21];
            mult_part_out12[186] <= P_5_4[5];
            mult_part_out12[187] <= P_7_2[20];
            mult_part_out12[188] <= P_6_3[14];
            mult_part_out12[189] <= P_3_5[18];
            mult_part_out12[190] <= P_6_3[16];
            mult_part_out12[191] <= P_0_7[23];
            mult_part_out12[192] <= P_0_7[24];
            mult_part_out12[193] <= P_3_5[22];
            mult_part_out12[194] <= P_10_1[0];
            mult_part_out12[195] <= P_0_7[27];
            mult_part_out12[196] <= P_2_6[18];
            mult_part_out12[197] <= P_7_3[6];
            mult_part_out12[198] <= P_9_1[21];
            mult_part_out12[199] <= P_10_1[5];
            mult_part_out12[200] <= P_0_8[8];
            mult_part_out12[201] <= P_11_0[14];
            mult_part_out12[202] <= P_4_5[14];
            mult_part_out12[203] <= P_5_4[22];
            mult_part_out12[204] <= P_7_2[37];
            mult_part_out12[205] <= P_1_7[20];
            mult_part_out12[206] <= P_2_7[4];
            mult_part_out12[207] <= P_5_5[2];
            mult_part_out12[208] <= P_7_3[17];
            mult_part_out12[209] <= P_5_5[4];
            mult_part_out12[210] <= P_6_3[36];
            mult_part_out12[211] <= P_3_6[16];
            mult_part_out12[212] <= P_4_6[0];
            mult_part_out12[213] <= P_6_3[39];
            mult_part_out12[214] <= P_2_7[12];
            mult_part_out12[215] <= P_7_4[0];
            mult_part_out12[216] <= P_2_6[38];
            mult_part_out12[217] <= P_5_4[36];
            mult_part_out12[218] <= P_9_2[17];
            mult_part_out12[219] <= P_2_7[17];
            mult_part_out12[220] <= P_0_8[28];
            mult_part_out12[221] <= P_2_7[19];
            mult_part_out12[222] <= P_10_2[4];
            mult_part_out12[223] <= P_1_7[38];
            mult_part_out12[224] <= P_3_6[29];
            mult_part_out12[225] <= P_11_1[14];
            mult_part_out12[226] <= P_11_1[15];
            mult_part_out12[227] <= P_9_2[26];
            mult_part_out12[228] <= P_5_5[23];
            mult_part_out12[229] <= P_0_8[37];
            mult_part_out12[230] <= P_10_2[12];
            mult_part_out12[231] <= P_9_3[6];
            mult_part_out12[232] <= P_3_7[13];
            mult_part_out12[233] <= P_3_6[38];
            mult_part_out12[234] <= P_2_8[8];
            mult_part_out12[235] <= P_13_0[14];
            mult_part_out12[236] <= P_1_9[3];
            mult_part_out12[237] <= P_9_2[36];
            mult_part_out12[238] <= P_3_7[19];
            mult_part_out12[239] <= P_11_2[4];
            mult_part_out12[240] <= P_1_8[31];
            mult_part_out12[241] <= P_14_0[3];
            mult_part_out12[242] <= P_4_6[30];
            mult_part_out12[243] <= P_1_9[10];
            mult_part_out12[244] <= P_2_8[18];
            mult_part_out12[245] <= P_11_2[10];
            mult_part_out12[246] <= P_13_1[1];
            mult_part_out12[247] <= P_10_2[29];
            mult_part_out12[248] <= P_4_6[36];
            mult_part_out12[249] <= P_7_4[34];
            mult_part_out12[250] <= P_14_0[12];
            mult_part_out12[251] <= P_4_6[39];
            mult_part_out12[252] <= P_5_6[23];
            mult_part_out12[253] <= P_8_4[21];
            mult_part_out12[254] <= P_12_2[2];
            mult_part_out12[255] <= P_4_7[19];
            mult_part_out12[256] <= P_10_2[38];
            mult_part_out12[257] <= P_2_9[7];
            mult_part_out12[258] <= P_1_10[1];
            mult_part_out12[259] <= P_5_7[6];
            mult_part_out12[260] <= P_3_8[17];
            mult_part_out12[261] <= P_8_5[5];
            mult_part_out12[262] <= P_4_7[26];
            mult_part_out12[263] <= P_2_9[13];
            mult_part_out12[264] <= P_11_2[29];
            mult_part_out12[265] <= P_8_5[9];
            mult_part_out12[266] <= P_2_9[16];
            mult_part_out12[267] <= P_11_3[8];
            mult_part_out12[268] <= P_10_3[26];
            mult_part_out12[269] <= P_4_7[33];
            mult_part_out12[270] <= P_12_2[18];
            mult_part_out12[271] <= P_9_4[22];
            mult_part_out12[272] <= P_10_4[6];
            mult_part_out12[273] <= P_11_3[14];
            mult_part_out12[274] <= P_3_9[7];
            mult_part_out12[275] <= P_12_2[23];
            mult_part_out12[276] <= P_5_7[23];
            mult_part_out12[277] <= P_7_5[38];
            mult_part_out12[278] <= P_2_10[4];
            mult_part_out12[279] <= P_9_4[30];
            mult_part_out12[280] <= P_10_4[14];
            mult_part_out12[281] <= P_6_6[35];
            mult_part_out12[282] <= P_5_8[5];
            mult_part_out12[283] <= P_2_10[9];
            mult_part_out12[284] <= P_12_3[8];
            mult_part_out12[285] <= P_5_7[32];
            mult_part_out12[286] <= P_12_2[34];
            mult_part_out12[287] <= P_6_7[17];
            mult_part_out12[288] <= P_8_6[8];
            mult_part_out12[289] <= P_7_6[26];
            mult_part_out12[290] <= P_2_9[40];
            mult_part_out12[291] <= P_3_9[24];
            mult_part_out12[292] <= P_7_7[5];
            mult_part_out12[293] <= P_3_10[2];
            mult_part_out12[294] <= P_14_1[32];
            mult_part_out12[295] <= P_14_1[33];
            mult_part_out12[296] <= P_13_3[3];
            mult_part_out12[297] <= P_11_3[38];
            mult_part_out12[298] <= P_14_1[36];
            mult_part_out12[299] <= P_6_8[5];
            mult_part_out12[300] <= P_10_5[10];
            mult_part_out12[301] <= P_13_2[32];
            mult_part_out12[302] <= P_4_9[18];
            mult_part_out12[303] <= P_9_5[30];
            mult_part_out12[304] <= P_15_2[1];
            mult_part_out12[305] <= P_13_2[36];
            mult_part_out12[306] <= P_3_10[15];
            mult_part_out12[307] <= P_7_7[20];
            mult_part_out12[308] <= P_12_3[32];
            mult_part_out12[309] <= P_10_5[19];
            mult_part_out12[310] <= P_12_3[34];
            mult_part_out12[311] <= P_11_5[4];
            mult_part_out12[312] <= P_9_6[15];
            mult_part_out12[313] <= P_9_6[16];
            mult_part_out12[314] <= P_4_9[30];
            mult_part_out12[315] <= P_11_4[32];
            mult_part_out12[316] <= P_5_8[39];
            mult_part_out12[317] <= P_4_9[33];
            mult_part_out12[318] <= P_8_6[38];
            mult_part_out12[319] <= P_7_7[32];
            mult_part_out12[320] <= P_13_3[27];
            mult_part_out12[321] <= P_4_10[13];
            mult_part_out12[322] <= P_14_2[36];
            mult_part_out12[323] <= P_9_6[26];
            mult_part_out12[324] <= P_14_3[14];
            mult_part_out12[325] <= P_11_5[18];
            mult_part_out12[326] <= P_12_5[2];
            mult_part_out12[327] <= P_10_6[13];
            mult_part_out12[328] <= P_10_5[38];
            mult_part_out12[329] <= P_8_7[25];
            mult_part_out12[330] <= P_7_8[19];
            mult_part_out12[331] <= P_6_8[37];
            mult_part_out12[332] <= P_9_6[35];
            mult_part_out12[333] <= P_5_10[8];
            mult_part_out12[334] <= P_7_8[23];
            mult_part_out12[335] <= P_14_4[1];
            mult_part_out12[336] <= P_12_5[12];
            mult_part_out12[337] <= P_13_4[20];
            mult_part_out12[338] <= P_8_7[34];
            mult_part_out12[339] <= P_14_3[29];
            mult_part_out12[340] <= P_7_8[29];
            mult_part_out12[341] <= P_11_5[34];
            mult_part_out12[342] <= P_13_5[1];
            mult_part_out12[343] <= P_11_5[36];
            mult_part_out12[344] <= P_9_7[23];
            mult_part_out12[345] <= P_10_7[7];
            mult_part_out12[346] <= P_13_5[5];
            mult_part_out12[347] <= P_11_5[40];
            mult_part_out12[348] <= P_6_10[6];
            mult_part_out12[349] <= P_13_4[32];
            mult_part_out12[350] <= P_10_6[36];
            mult_part_out12[351] <= P_6_10[9];
            mult_part_out12[352] <= P_13_4[35];
            mult_part_out12[353] <= P_10_7[15];
            mult_part_out12[354] <= P_10_7[16];
            mult_part_out12[355] <= P_8_9[3];
            mult_part_out12[356] <= P_9_7[35];
            mult_part_out12[357] <= P_6_10[15];
            mult_part_out12[358] <= P_7_9[23];
            mult_part_out12[359] <= P_15_4[8];
            mult_part_out12[360] <= P_12_6[12];
            mult_part_out12[361] <= P_11_7[6];
            mult_part_out12[362] <= P_8_9[10];
            mult_part_out12[363] <= P_14_5[5];
            mult_part_out12[364] <= P_14_4[30];
            mult_part_out12[365] <= P_8_9[13];
            mult_part_out12[366] <= P_15_4[15];
            mult_part_out12[367] <= P_12_6[19];
            mult_part_out12[368] <= P_11_7[13];
            mult_part_out12[369] <= P_15_4[18];
            mult_part_out12[370] <= P_7_9[35];
            mult_part_out12[371] <= P_7_10[12];
            mult_part_out12[372] <= P_14_5[14];
            mult_part_out12[373] <= P_13_5[32];
            mult_part_out12[374] <= P_14_4[40];
            mult_part_out12[375] <= P_7_9[40];
            mult_part_out12[376] <= P_12_6[28];
            mult_part_out12[377] <= P_9_9[8];
            mult_part_out12[378] <= P_15_5[3];
            mult_part_out12[379] <= P_10_8[17];
            mult_part_out12[380] <= P_13_5[39];
            mult_part_out12[381] <= P_13_6[16];
            mult_part_out12[382] <= P_7_10[23];
            mult_part_out12[383] <= P_7_10[24];
            mult_part_out12[384] <= P_8_10[8];
            mult_part_out12[385] <= P_13_6[20];
            mult_part_out12[386] <= P_8_10[10];
            mult_part_out12[387] <= P_10_9[1];
            mult_part_out12[388] <= P_14_6[6];
            mult_part_out12[389] <= P_7_10[30];
            mult_part_out12[390] <= P_11_8[11];
            mult_part_out12[391] <= P_10_9[5];
            mult_part_out12[392] <= P_11_8[13];
            mult_part_out12[393] <= P_14_6[11];
            mult_part_out12[394] <= P_13_6[29];
            mult_part_out12[395] <= P_9_9[26];
            mult_part_out12[396] <= P_9_9[27];
            mult_part_out12[397] <= P_11_8[18];
            mult_part_out12[398] <= P_12_7[26];
            mult_part_out12[399] <= P_9_9[30];

            mult_part_out13[136] <= P_4_2[20];
            mult_part_out13[137] <= P_1_4[24];
            mult_part_out13[138] <= P_0_5[18];
            mult_part_out13[139] <= P_3_3[16];
            mult_part_out13[140] <= P_2_4[10];
            mult_part_out13[141] <= P_4_3[1];
            mult_part_out13[142] <= P_4_2[26];
            mult_part_out13[143] <= P_1_4[30];
            mult_part_out13[144] <= P_2_3[38];
            mult_part_out13[145] <= P_3_3[22];
            mult_part_out13[146] <= P_5_2[13];
            mult_part_out13[147] <= P_1_4[34];
            mult_part_out13[148] <= P_3_3[25];
            mult_part_out13[149] <= P_3_3[26];
            mult_part_out13[150] <= P_3_4[3];
            mult_part_out13[151] <= P_3_3[28];
            mult_part_out13[152] <= P_8_0[16];
            mult_part_out13[153] <= P_7_0[34];
            mult_part_out13[154] <= P_0_6[10];
            mult_part_out13[155] <= P_7_1[12];
            mult_part_out13[156] <= P_9_0[3];
            mult_part_out13[157] <= P_3_3[34];
            mult_part_out13[158] <= P_0_5[38];
            mult_part_out13[159] <= P_5_3[2];
            mult_part_out13[160] <= P_0_6[16];
            mult_part_out13[161] <= P_0_6[17];
            mult_part_out13[162] <= P_0_6[18];
            mult_part_out13[163] <= P_5_2[30];
            mult_part_out13[164] <= P_1_6[3];
            mult_part_out13[165] <= P_6_1[39];
            mult_part_out13[166] <= P_4_3[26];
            mult_part_out13[167] <= P_7_2[0];
            mult_part_out13[168] <= P_9_0[15];
            mult_part_out13[169] <= P_5_3[12];
            mult_part_out13[170] <= P_8_1[10];
            mult_part_out13[171] <= P_8_0[35];
            mult_part_out13[172] <= P_3_5[1];
            mult_part_out13[173] <= P_7_1[30];
            mult_part_out13[174] <= P_1_5[37];
            mult_part_out13[175] <= P_3_5[4];
            mult_part_out13[176] <= P_9_0[23];
            mult_part_out13[177] <= P_9_0[24];
            mult_part_out13[178] <= P_2_6[0];
            mult_part_out13[179] <= P_3_4[32];
            mult_part_out13[180] <= P_3_4[33];
            mult_part_out13[181] <= P_5_3[24];
            mult_part_out13[182] <= P_7_2[15];
            mult_part_out13[183] <= P_2_5[29];
            mult_part_out13[184] <= P_2_5[30];
            mult_part_out13[185] <= P_5_4[4];
            mult_part_out13[186] <= P_8_2[2];
            mult_part_out13[187] <= P_4_4[23];
            mult_part_out13[188] <= P_8_1[28];
            mult_part_out13[189] <= P_4_4[25];
            mult_part_out13[190] <= P_6_2[40];
            mult_part_out13[191] <= P_10_0[21];
            mult_part_out13[192] <= P_4_4[28];
            mult_part_out13[193] <= P_0_7[25];
            mult_part_out13[194] <= P_5_4[13];
            mult_part_out13[195] <= P_4_4[31];
            mult_part_out13[196] <= P_4_4[32];
            mult_part_out13[197] <= P_8_2[13];
            mult_part_out13[198] <= P_2_6[20];
            mult_part_out13[199] <= P_4_5[11];
            mult_part_out13[200] <= P_1_7[15];
            mult_part_out13[201] <= P_0_7[33];
            mult_part_out13[202] <= P_0_8[10];
            mult_part_out13[203] <= P_10_0[33];
            mult_part_out13[204] <= P_2_6[26];
            mult_part_out13[205] <= P_8_2[21];
            mult_part_out13[206] <= P_0_8[14];
            mult_part_out13[207] <= P_6_3[33];
            mult_part_out13[208] <= P_3_5[37];
            mult_part_out13[209] <= P_3_5[38];
            mult_part_out13[210] <= P_6_4[12];
            mult_part_out13[211] <= P_8_2[27];
            mult_part_out13[212] <= P_8_2[28];
            mult_part_out13[213] <= P_4_5[25];
            mult_part_out13[214] <= P_4_6[2];
            mult_part_out13[215] <= P_1_7[30];
            mult_part_out13[216] <= P_11_0[29];
            mult_part_out13[217] <= P_2_6[39];
            mult_part_out13[218] <= P_4_5[30];
            mult_part_out13[219] <= P_8_2[35];
            mult_part_out13[220] <= P_3_7[1];
            mult_part_out13[221] <= P_9_2[20];
            mult_part_out13[222] <= P_3_7[3];
            mult_part_out13[223] <= P_2_7[21];
            mult_part_out13[224] <= P_6_4[26];
            mult_part_out13[225] <= P_9_3[0];
            mult_part_out13[226] <= P_11_0[39];
            mult_part_out13[227] <= P_7_3[36];
            mult_part_out13[228] <= P_13_0[7];
            mult_part_out13[229] <= P_8_3[21];
            mult_part_out13[230] <= P_2_8[4];
            mult_part_out13[231] <= P_12_1[3];
            mult_part_out13[232] <= P_0_8[40];
            mult_part_out13[233] <= P_8_4[1];
            mult_part_out13[234] <= P_5_5[29];
            mult_part_out13[235] <= P_6_4[37];
            mult_part_out13[236] <= P_2_8[10];
            mult_part_out13[237] <= P_11_1[26];
            mult_part_out13[238] <= P_5_5[33];
            mult_part_out13[239] <= P_9_2[38];
            mult_part_out13[240] <= P_6_5[18];
            mult_part_out13[241] <= P_6_5[19];
            mult_part_out13[242] <= P_5_5[37];
            mult_part_out13[243] <= P_7_5[4];
            mult_part_out13[244] <= P_0_10[4];
            mult_part_out13[245] <= P_0_9[29];
            mult_part_out13[246] <= P_7_4[31];
            mult_part_out13[247] <= P_14_0[9];
            mult_part_out13[248] <= P_10_2[30];
            mult_part_out13[249] <= P_10_3[7];
            mult_part_out13[250] <= P_10_3[8];
            mult_part_out13[251] <= P_10_2[33];
            mult_part_out13[252] <= P_9_3[27];
            mult_part_out13[253] <= P_3_8[10];
            mult_part_out13[254] <= P_14_0[16];
            mult_part_out13[255] <= P_2_8[29];
            mult_part_out13[256] <= P_2_8[30];
            mult_part_out13[257] <= P_11_2[22];
            mult_part_out13[258] <= P_8_4[26];
            mult_part_out13[259] <= P_8_5[3];
            mult_part_out13[260] <= P_4_7[24];
            mult_part_out13[261] <= P_4_8[1];
            mult_part_out13[262] <= P_6_6[16];
            mult_part_out13[263] <= P_11_2[28];
            mult_part_out13[264] <= P_9_3[39];
            mult_part_out13[265] <= P_3_8[22];
            mult_part_out13[266] <= P_9_4[17];
            mult_part_out13[267] <= P_5_7[14];
            mult_part_out13[268] <= P_8_5[12];
            mult_part_out13[269] <= P_5_6[40];
            mult_part_out13[270] <= P_11_2[35];
            mult_part_out13[271] <= P_5_7[18];
            mult_part_out13[272] <= P_14_0[34];
            mult_part_out13[273] <= P_9_5[0];
            mult_part_out13[274] <= P_13_1[29];
            mult_part_out13[275] <= P_14_0[37];
            mult_part_out13[276] <= P_8_5[20];
            mult_part_out13[277] <= P_2_10[3];
            mult_part_out13[278] <= P_15_0[23];
            mult_part_out13[279] <= P_10_4[13];
            mult_part_out13[280] <= P_12_3[4];
            mult_part_out13[281] <= P_3_9[14];
            mult_part_out13[282] <= P_3_8[39];
            mult_part_out13[283] <= P_3_9[16];
            mult_part_out13[284] <= P_7_6[21];
            mult_part_out13[285] <= P_9_5[12];
            mult_part_out13[286] <= P_3_9[19];
            mult_part_out13[287] <= P_2_9[37];
            mult_part_out13[288] <= P_14_2[2];
            mult_part_out13[289] <= P_4_9[5];
            mult_part_out13[290] <= P_5_8[13];
            mult_part_out13[291] <= P_15_1[12];
            mult_part_out13[292] <= P_14_1[30];
            mult_part_out13[293] <= P_4_9[9];
            mult_part_out13[294] <= P_11_4[11];
            mult_part_out13[295] <= P_5_8[18];
            mult_part_out13[296] <= P_8_5[40];
            mult_part_out13[297] <= P_15_1[18];
            mult_part_out13[298] <= P_8_6[18];
            mult_part_out13[299] <= P_13_3[6];
            mult_part_out13[300] <= P_6_7[30];
            mult_part_out13[301] <= P_5_9[0];
            mult_part_out13[302] <= P_6_7[32];
            mult_part_out13[303] <= P_13_3[10];
            mult_part_out13[304] <= P_12_4[4];
            mult_part_out13[305] <= P_4_9[21];
            mult_part_out13[306] <= P_5_8[29];
            mult_part_out13[307] <= P_5_8[30];
            mult_part_out13[308] <= P_5_8[31];
            mult_part_out13[309] <= P_7_7[22];
            mult_part_out13[310] <= P_12_4[10];
            mult_part_out13[311] <= P_15_2[8];
            mult_part_out13[312] <= P_8_7[8];
            mult_part_out13[313] <= P_9_5[40];
            mult_part_out13[314] <= P_7_7[27];
            mult_part_out13[315] <= P_13_3[22];
            mult_part_out13[316] <= P_15_2[13];
            mult_part_out13[317] <= P_6_8[23];
            mult_part_out13[318] <= P_7_8[7];
            mult_part_out13[319] <= P_10_5[29];
            mult_part_out13[320] <= P_13_4[3];
            mult_part_out13[321] <= P_7_7[34];
            mult_part_out13[322] <= P_11_4[39];
            mult_part_out13[323] <= P_7_7[36];
            mult_part_out13[324] <= P_4_9[40];
            mult_part_out13[325] <= P_10_6[11];
            mult_part_out13[326] <= P_13_4[9];
            mult_part_out13[327] <= P_6_8[33];
            mult_part_out13[328] <= P_6_9[10];
            mult_part_out13[329] <= P_7_8[18];
            mult_part_out13[330] <= P_12_4[30];
            mult_part_out13[331] <= P_6_9[13];
            mult_part_out13[332] <= P_15_3[5];
            mult_part_out13[333] <= P_15_3[6];
            mult_part_out13[334] <= P_11_5[27];
            mult_part_out13[335] <= P_7_8[24];
            mult_part_out13[336] <= P_9_7[15];
            mult_part_out13[337] <= P_7_8[26];
            mult_part_out13[338] <= P_13_4[21];
            mult_part_out13[339] <= P_7_9[4];
            mult_part_out13[340] <= P_8_7[36];
            mult_part_out13[341] <= P_14_3[31];
            mult_part_out13[342] <= P_7_8[31];
            mult_part_out13[343] <= P_7_8[32];
            mult_part_out13[344] <= P_8_8[16];
            mult_part_out13[345] <= P_14_4[11];
            mult_part_out13[346] <= P_6_9[28];
            mult_part_out13[347] <= P_15_3[20];
            mult_part_out13[348] <= P_12_5[24];
            mult_part_out13[349] <= P_10_6[35];
            mult_part_out13[350] <= P_11_6[19];
            mult_part_out13[351] <= P_12_5[27];
            mult_part_out13[352] <= P_8_8[24];
            mult_part_out13[353] <= P_8_9[1];
            mult_part_out13[354] <= P_10_6[40];
            mult_part_out13[355] <= P_8_8[27];
            mult_part_out13[356] <= P_11_7[1];
            mult_part_out13[357] <= P_15_4[6];
            mult_part_out13[358] <= P_6_10[16];
            mult_part_out13[359] <= P_7_9[24];
            mult_part_out13[360] <= P_7_9[25];
            mult_part_out13[361] <= P_8_8[33];
            mult_part_out13[362] <= P_7_9[27];
            mult_part_out13[363] <= P_12_5[39];
            mult_part_out13[364] <= P_14_5[6];
            mult_part_out13[365] <= P_15_4[14];
            mult_part_out13[366] <= P_10_7[28];
            mult_part_out13[367] <= P_7_10[8];
            mult_part_out13[368] <= P_8_9[16];
            mult_part_out13[369] <= P_10_7[31];
            mult_part_out13[370] <= P_14_4[36];
            mult_part_out13[371] <= P_11_6[40];
            mult_part_out13[372] <= P_6_10[30];
            mult_part_out13[373] <= P_10_8[11];
            mult_part_out13[374] <= P_7_9[39];
            mult_part_out13[375] <= P_13_5[34];
            mult_part_out13[376] <= P_8_10[0];
            mult_part_out13[377] <= P_8_9[25];
            mult_part_out13[378] <= P_12_7[6];
            mult_part_out13[379] <= P_11_8[0];
            mult_part_out13[380] <= P_12_7[8];
            mult_part_out13[381] <= P_8_10[5];
            mult_part_out13[382] <= P_14_6[0];
            mult_part_out13[383] <= P_9_9[14];
            mult_part_out13[384] <= P_11_8[5];
            mult_part_out13[385] <= P_11_7[30];
            mult_part_out13[386] <= P_11_8[7];
            mult_part_out13[387] <= P_9_9[18];
            mult_part_out13[388] <= P_8_10[12];
            mult_part_out13[389] <= P_8_9[37];
            mult_part_out13[390] <= P_14_6[8];
            mult_part_out13[391] <= P_15_5[16];

            mult_part_out14[144] <= P_6_1[18];
            mult_part_out14[145] <= P_5_1[36];
            mult_part_out14[146] <= P_2_3[40];
            mult_part_out14[147] <= P_7_0[28];
            mult_part_out14[148] <= P_0_5[28];
            mult_part_out14[149] <= P_0_5[29];
            mult_part_out14[150] <= P_6_2[0];
            mult_part_out14[151] <= P_0_5[31];
            mult_part_out14[152] <= P_0_6[8];
            mult_part_out14[153] <= P_1_5[16];
            mult_part_out14[154] <= P_6_2[4];
            mult_part_out14[155] <= P_4_3[15];
            mult_part_out14[156] <= P_4_2[40];
            mult_part_out14[157] <= P_7_0[38];
            mult_part_out14[158] <= P_6_1[32];
            mult_part_out14[159] <= P_2_4[29];
            mult_part_out14[160] <= P_2_5[6];
            mult_part_out14[161] <= P_5_2[28];
            mult_part_out14[162] <= P_7_1[19];
            mult_part_out14[163] <= P_3_4[16];
            mult_part_out14[164] <= P_3_4[17];
            mult_part_out14[165] <= P_0_6[21];
            mult_part_out14[166] <= P_5_3[9];
            mult_part_out14[167] <= P_1_6[6];
            mult_part_out14[168] <= P_4_4[4];
            mult_part_out14[169] <= P_2_5[15];
            mult_part_out14[170] <= P_7_2[3];
            mult_part_out14[171] <= P_9_0[18];
            mult_part_out14[172] <= P_6_2[22];
            mult_part_out14[173] <= P_7_2[6];
            mult_part_out14[174] <= P_8_1[14];
            mult_part_out14[175] <= P_4_4[11];
            mult_part_out14[176] <= P_6_2[26];
            mult_part_out14[177] <= P_1_6[16];
            mult_part_out14[178] <= P_6_2[28];
            mult_part_out14[179] <= P_7_2[12];
            mult_part_out14[180] <= P_6_2[30];
            mult_part_out14[181] <= P_3_5[10];
            mult_part_out14[182] <= P_2_5[28];
            mult_part_out14[183] <= P_2_6[5];
            mult_part_out14[184] <= P_0_7[16];
            mult_part_out14[185] <= P_2_5[31];
            mult_part_out14[186] <= P_1_6[25];
            mult_part_out14[187] <= P_3_5[16];
            mult_part_out14[188] <= P_2_6[10];
            mult_part_out14[189] <= P_10_0[19];
            mult_part_out14[190] <= P_8_1[30];
            mult_part_out14[191] <= P_8_2[7];
            mult_part_out14[192] <= P_8_1[32];
            mult_part_out14[193] <= P_1_6[32];
            mult_part_out14[194] <= P_5_3[37];
            mult_part_out14[195] <= P_4_5[7];
            mult_part_out14[196] <= P_0_8[4];
            mult_part_out14[197] <= P_11_0[10];
            mult_part_out14[198] <= P_4_4[34];
            mult_part_out14[199] <= P_5_4[18];
            mult_part_out14[200] <= P_7_2[33];
            mult_part_out14[201] <= P_5_4[20];
            mult_part_out14[202] <= P_9_1[25];
            mult_part_out14[203] <= P_9_2[2];
            mult_part_out14[204] <= P_7_3[13];
            mult_part_out14[205] <= P_5_4[24];
            mult_part_out14[206] <= P_12_0[2];
            mult_part_out14[207] <= P_10_0[37];
            mult_part_out14[208] <= P_2_6[30];
            mult_part_out14[209] <= P_6_4[11];
            mult_part_out14[210] <= P_11_0[23];
            mult_part_out14[211] <= P_9_1[34];
            mult_part_out14[212] <= P_3_6[17];
            mult_part_out14[213] <= P_9_1[36];
            mult_part_out14[214] <= P_5_5[9];
            mult_part_out14[215] <= P_6_4[17];
            mult_part_out14[216] <= P_4_5[28];
            mult_part_out14[217] <= P_1_8[8];
            mult_part_out14[218] <= P_5_4[37];
            mult_part_out14[219] <= P_6_4[21];
            mult_part_out14[220] <= P_5_4[39];
            mult_part_out14[221] <= P_11_1[10];
            mult_part_out14[222] <= P_8_3[14];
            mult_part_out14[223] <= P_9_2[22];
            mult_part_out14[224] <= P_1_7[39];
            mult_part_out14[225] <= P_1_7[40];
            mult_part_out14[226] <= P_13_0[5];
            mult_part_out14[227] <= P_3_7[8];
            mult_part_out14[228] <= P_0_9[12];
            mult_part_out14[229] <= P_5_5[24];
            mult_part_out14[230] <= P_2_7[28];
            mult_part_out14[231] <= P_8_3[23];
            mult_part_out14[232] <= P_10_1[38];
            mult_part_out14[233] <= P_10_1[39];
            mult_part_out14[234] <= P_6_4[36];
            mult_part_out14[235] <= P_1_8[26];
            mult_part_out14[236] <= P_8_4[4];
            mult_part_out14[237] <= P_10_2[19];
            mult_part_out14[238] <= P_4_6[26];
            mult_part_out14[239] <= P_12_0[35];
            mult_part_out14[240] <= P_14_0[2];
            mult_part_out14[241] <= P_1_9[8];
            mult_part_out14[242] <= P_8_4[10];
            mult_part_out14[243] <= P_10_3[1];
            mult_part_out14[244] <= P_7_4[29];
            mult_part_out14[245] <= P_7_5[6];
            mult_part_out14[246] <= P_3_8[3];
            mult_part_out14[247] <= P_4_6[35];
            mult_part_out14[248] <= P_7_5[9];
            mult_part_out14[249] <= P_4_6[37];
            mult_part_out14[250] <= P_10_2[32];
            mult_part_out14[251] <= P_5_6[22];
            mult_part_out14[252] <= P_12_2[0];
            mult_part_out14[253] <= P_9_4[4];
            mult_part_out14[254] <= P_2_9[4];
            mult_part_out14[255] <= P_6_6[9];
            mult_part_out14[256] <= P_3_7[37];
            mult_part_out14[257] <= P_13_1[12];
            mult_part_out14[258] <= P_12_1[30];
            mult_part_out14[259] <= P_5_6[30];
            mult_part_out14[260] <= P_1_9[27];
            mult_part_out14[261] <= P_2_8[35];
            mult_part_out14[262] <= P_7_5[23];
            mult_part_out14[263] <= P_1_10[6];
            mult_part_out14[264] <= P_4_7[28];
            mult_part_out14[265] <= P_7_5[26];
            mult_part_out14[266] <= P_13_1[21];
            mult_part_out14[267] <= P_12_2[15];
            mult_part_out14[268] <= P_9_4[19];
            mult_part_out14[269] <= P_5_7[16];
            mult_part_out14[270] <= P_1_9[37];
            mult_part_out14[271] <= P_15_0[16];
            mult_part_out14[272] <= P_3_8[29];
            mult_part_out14[273] <= P_1_10[16];
            mult_part_out14[274] <= P_6_6[28];
            mult_part_out14[275] <= P_5_7[22];
            mult_part_out14[276] <= P_1_10[19];
            mult_part_out14[277] <= P_8_5[21];
            mult_part_out14[278] <= P_3_9[11];
            mult_part_out14[279] <= P_3_9[12];
            mult_part_out14[280] <= P_6_6[34];
            mult_part_out14[281] <= P_12_2[29];
            mult_part_out14[282] <= P_1_10[25];
            mult_part_out14[283] <= P_13_2[14];
            mult_part_out14[284] <= P_6_6[38];
            mult_part_out14[285] <= P_2_10[11];
            mult_part_out14[286] <= P_2_10[12];
            mult_part_out14[287] <= P_2_10[13];
            mult_part_out14[288] <= P_12_2[36];
            mult_part_out14[289] <= P_8_6[9];
            mult_part_out14[290] <= P_14_2[4];
            mult_part_out14[291] <= P_14_1[29];
            mult_part_out14[292] <= P_4_9[8];
            mult_part_out14[293] <= P_10_5[3];
            mult_part_out14[294] <= P_5_8[17];
            mult_part_out14[295] <= P_4_9[11];
            mult_part_out14[296] <= P_10_5[6];
            mult_part_out14[297] <= P_11_4[14];
            mult_part_out14[298] <= P_14_2[12];
            mult_part_out14[299] <= P_11_4[16];
            mult_part_out14[300] <= P_15_1[21];
            mult_part_out14[301] <= P_2_10[27];
            mult_part_out14[302] <= P_7_6[39];
            mult_part_out14[303] <= P_5_9[2];
            mult_part_out14[304] <= P_9_6[7];
            mult_part_out14[305] <= P_5_8[28];
            mult_part_out14[306] <= P_6_7[36];
            mult_part_out14[307] <= P_12_4[7];
            mult_part_out14[308] <= P_13_3[15];
            mult_part_out14[309] <= P_5_8[32];
            mult_part_out14[310] <= P_15_2[7];
            mult_part_out14[311] <= P_8_7[7];
            mult_part_out14[312] <= P_4_10[4];
            mult_part_out14[313] <= P_11_5[6];
            mult_part_out14[314] <= P_8_7[10];
            mult_part_out14[315] <= P_5_8[38];
            mult_part_out14[316] <= P_7_8[5];
            mult_part_out14[317] <= P_14_3[7];
            mult_part_out14[318] <= P_14_2[32];
            mult_part_out14[319] <= P_8_7[15];
            mult_part_out14[320] <= P_11_4[37];
            mult_part_out14[321] <= P_9_7[0];
            mult_part_out14[322] <= P_4_10[14];
            mult_part_out14[323] <= P_15_2[20];
            mult_part_out14[324] <= P_9_7[3];
            mult_part_out14[325] <= P_14_3[15];
            mult_part_out14[326] <= P_8_7[22];
            mult_part_out14[327] <= P_4_10[19];
            mult_part_out14[328] <= P_4_10[20];
            mult_part_out14[329] <= P_13_4[12];
            mult_part_out14[330] <= P_13_4[13];
            mult_part_out14[331] <= P_8_8[3];
            mult_part_out14[332] <= P_12_5[8];
            mult_part_out14[333] <= P_5_9[32];
            mult_part_out14[334] <= P_15_3[7];
            mult_part_out14[335] <= P_11_5[28];
            mult_part_out14[336] <= P_10_6[22];
            mult_part_out14[337] <= P_11_6[6];
            mult_part_out14[338] <= P_12_5[14];
            mult_part_out14[339] <= P_13_4[22];
            mult_part_out14[340] <= P_5_9[39];
            mult_part_out14[341] <= P_13_5[0];
            mult_part_out14[342] <= P_10_6[28];
            mult_part_out14[343] <= P_10_7[5];
            mult_part_out14[344] <= P_14_3[34];
            mult_part_out14[345] <= P_15_3[18];
            mult_part_out14[346] <= P_8_8[18];
            mult_part_out14[347] <= P_7_9[12];
            mult_part_out14[348] <= P_13_5[7];
            mult_part_out14[349] <= P_11_6[18];
            mult_part_out14[350] <= P_9_8[5];
            mult_part_out14[351] <= P_15_4[0];
            mult_part_out14[352] <= P_5_10[27];
            mult_part_out14[353] <= P_13_5[12];
            mult_part_out14[354] <= P_9_7[33];
            mult_part_out14[355] <= P_11_6[24];
            mult_part_out14[356] <= P_7_9[21];
            mult_part_out14[357] <= P_13_4[40];
            mult_part_out14[358] <= P_8_9[6];
            mult_part_out14[359] <= P_12_6[11];
            mult_part_out14[360] <= P_13_5[19];
            mult_part_out14[361] <= P_12_5[37];
            mult_part_out14[362] <= P_14_4[28];
            mult_part_out14[363] <= P_7_10[4];
            mult_part_out14[364] <= P_8_9[12];
            mult_part_out14[365] <= P_7_10[6];
            mult_part_out14[366] <= P_11_6[35];
            mult_part_out14[367] <= P_10_8[5];
            mult_part_out14[368] <= P_10_8[6];
            mult_part_out14[369] <= P_8_9[17];
            mult_part_out14[370] <= P_10_7[32];
            mult_part_out14[371] <= P_14_5[13];
            mult_part_out14[372] <= P_10_7[34];
            mult_part_out14[373] <= P_6_10[31];
            mult_part_out14[374] <= P_14_5[16];
            mult_part_out14[375] <= P_15_5[0];

            mult_part_out15[153] <= P_6_2[3];
            mult_part_out15[154] <= P_7_0[35];
            mult_part_out15[155] <= P_6_2[5];
            mult_part_out15[156] <= P_2_5[2];
            mult_part_out15[157] <= P_8_0[21];
            mult_part_out15[158] <= P_1_5[21];
            mult_part_out15[159] <= P_3_4[12];
            mult_part_out15[160] <= P_7_1[17];
            mult_part_out15[161] <= P_2_5[7];
            mult_part_out15[162] <= P_1_5[25];
            mult_part_out15[163] <= P_7_1[20];
            mult_part_out15[164] <= P_2_5[10];
            mult_part_out15[165] <= P_1_5[28];
            mult_part_out15[166] <= P_2_4[36];
            mult_part_out15[167] <= P_5_2[34];
            mult_part_out15[168] <= P_1_6[7];
            mult_part_out15[169] <= P_3_4[22];
            mult_part_out15[170] <= P_10_0[0];
            mult_part_out15[171] <= P_10_0[1];
            mult_part_out15[172] <= P_1_6[11];
            mult_part_out15[173] <= P_3_5[2];
            mult_part_out15[174] <= P_8_0[38];
            mult_part_out15[175] <= P_0_6[31];
            mult_part_out15[176] <= P_8_0[40];
            mult_part_out15[177] <= P_5_3[20];
            mult_part_out15[178] <= P_2_5[24];
            mult_part_out15[179] <= P_5_3[22];
            mult_part_out15[180] <= P_6_3[6];
            mult_part_out15[181] <= P_3_4[34];
            mult_part_out15[182] <= P_10_0[12];
            mult_part_out15[183] <= P_0_6[39];
            mult_part_out15[184] <= P_6_2[34];
            mult_part_out15[185] <= P_2_6[7];
            mult_part_out15[186] <= P_0_7[18];
            mult_part_out15[187] <= P_8_1[27];
            mult_part_out15[188] <= P_4_5[0];
            mult_part_out15[189] <= P_1_6[28];
            mult_part_out15[190] <= P_8_2[6];
            mult_part_out15[191] <= P_5_3[34];
            mult_part_out15[192] <= P_11_0[5];
            mult_part_out15[193] <= P_4_4[29];
            mult_part_out15[194] <= P_4_5[6];
            mult_part_out15[195] <= P_1_6[34];
            mult_part_out15[196] <= P_10_0[26];
            mult_part_out15[197] <= P_5_4[16];
            mult_part_out15[198] <= P_0_8[6];
            mult_part_out15[199] <= P_8_2[15];
            mult_part_out15[200] <= P_11_0[13];
            mult_part_out15[201] <= P_0_8[9];
            mult_part_out15[202] <= P_4_4[38];
            mult_part_out15[203] <= P_0_8[11];
            mult_part_out15[204] <= P_9_1[27];
            mult_part_out15[205] <= P_0_7[37];
            mult_part_out15[206] <= P_3_5[35];
            mult_part_out15[207] <= P_0_7[39];
            mult_part_out15[208] <= P_9_1[31];
            mult_part_out15[209] <= P_10_1[15];
            mult_part_out15[210] <= P_3_6[15];
            mult_part_out15[211] <= P_6_3[37];
            mult_part_out15[212] <= P_12_0[8];
            mult_part_out15[213] <= P_7_3[22];
            mult_part_out15[214] <= P_2_6[36];
            mult_part_out15[215] <= P_7_3[24];
            mult_part_out15[216] <= P_12_0[12];
            mult_part_out15[217] <= P_9_2[16];
            mult_part_out15[218] <= P_8_2[34];
            mult_part_out15[219] <= P_10_1[25];
            mult_part_out15[220] <= P_9_2[19];
            mult_part_out15[221] <= P_5_5[16];
            mult_part_out15[222] <= P_0_9[6];
            mult_part_out15[223] <= P_7_3[32];
            mult_part_out15[224] <= P_10_2[6];
            mult_part_out15[225] <= P_7_4[10];
            mult_part_out15[226] <= P_8_3[18];
            mult_part_out15[227] <= P_9_3[2];
            mult_part_out15[228] <= P_4_6[16];
            mult_part_out15[229] <= P_3_7[10];
            mult_part_out15[230] <= P_10_1[36];
            mult_part_out15[231] <= P_1_8[22];
            mult_part_out15[232] <= P_8_4[0];
            mult_part_out15[233] <= P_8_3[25];
            mult_part_out15[234] <= P_9_2[33];
            mult_part_out15[235] <= P_8_4[3];
            mult_part_out15[236] <= P_8_3[28];
            mult_part_out15[237] <= P_1_9[4];
            mult_part_out15[238] <= P_11_1[27];
            mult_part_out15[239] <= P_9_3[14];
            mult_part_out15[240] <= P_0_9[24];
            mult_part_out15[241] <= P_1_8[32];
            mult_part_out15[242] <= P_4_7[6];
            mult_part_out15[243] <= P_8_4[11];
            mult_part_out15[244] <= P_5_5[39];
            mult_part_out15[245] <= P_4_7[9];
            mult_part_out15[246] <= P_2_8[20];
            mult_part_out15[247] <= P_5_6[18];
            mult_part_out15[248] <= P_10_3[6];
            mult_part_out15[249] <= P_7_5[10];
            mult_part_out15[250] <= P_7_4[35];
            mult_part_out15[251] <= P_3_8[8];
            mult_part_out15[252] <= P_1_9[19];
            mult_part_out15[253] <= P_6_6[7];
            mult_part_out15[254] <= P_1_9[21];
            mult_part_out15[255] <= P_3_8[12];
            mult_part_out15[256] <= P_8_4[24];
            mult_part_out15[257] <= P_5_7[4];
            mult_part_out15[258] <= P_3_7[39];
            mult_part_out15[259] <= P_11_3[0];
            mult_part_out15[260] <= P_7_5[21];
            mult_part_out15[261] <= P_12_2[9];
            mult_part_out15[262] <= P_9_4[13];
            mult_part_out15[263] <= P_8_5[7];
            mult_part_out15[264] <= P_2_9[14];
            mult_part_out15[265] <= P_7_6[2];
            mult_part_out15[266] <= P_11_2[31];
            mult_part_out15[267] <= P_3_8[24];
            mult_part_out15[268] <= P_6_6[22];
            mult_part_out15[269] <= P_12_2[17];
            mult_part_out15[270] <= P_13_2[1];
            mult_part_out15[271] <= P_7_6[8];
            mult_part_out15[272] <= P_6_6[26];
            mult_part_out15[273] <= P_7_6[10];
            mult_part_out15[274] <= P_10_3[32];
            mult_part_out15[275] <= P_8_5[19];
            mult_part_out15[276] <= P_6_7[6];
            mult_part_out15[277] <= P_13_2[8];
            mult_part_out15[278] <= P_10_4[12];
            mult_part_out15[279] <= P_12_3[3];
            mult_part_out15[280] <= P_9_5[7];
            mult_part_out15[281] <= P_10_3[39];
            mult_part_out15[282] <= P_3_9[15];
            mult_part_out15[283] <= P_9_4[34];
            mult_part_out15[284] <= P_4_8[24];
            mult_part_out15[285] <= P_13_2[16];
            mult_part_out15[286] <= P_12_3[10];
            mult_part_out15[287] <= P_4_9[3];
            mult_part_out15[288] <= P_2_10[14];
            mult_part_out15[289] <= P_4_8[29];
            mult_part_out15[290] <= P_8_6[10];
            mult_part_out15[291] <= P_4_9[7];
            mult_part_out15[292] <= P_10_4[26];
            mult_part_out15[293] <= P_11_4[10];
            mult_part_out15[294] <= P_12_3[18];
            mult_part_out15[295] <= P_6_8[1];
            mult_part_out15[296] <= P_14_1[34];
            mult_part_out15[297] <= P_5_8[20];
            mult_part_out15[298] <= P_15_1[19];
            mult_part_out15[299] <= P_14_1[37];
            mult_part_out15[300] <= P_2_10[26];
            mult_part_out15[301] <= P_8_6[21];
            mult_part_out15[302] <= P_14_1[40];
            mult_part_out15[303] <= P_5_8[26];
            mult_part_out15[304] <= P_10_5[14];
            mult_part_out15[305] <= P_12_4[5];
            mult_part_out15[306] <= P_6_8[12];
            mult_part_out15[307] <= P_6_8[13];
            mult_part_out15[308] <= P_14_2[22];
            mult_part_out15[309] <= P_5_9[8];
            mult_part_out15[310] <= P_9_5[37];
            mult_part_out15[311] <= P_10_5[21];
            mult_part_out15[312] <= P_14_2[26];
            mult_part_out15[313] <= P_3_10[22];
            mult_part_out15[314] <= P_7_8[3];
            mult_part_out15[315] <= P_15_2[12];
            mult_part_out15[316] <= P_3_10[25];
            mult_part_out15[317] <= P_8_7[13];
            mult_part_out15[318] <= P_15_2[15];
            mult_part_out15[319] <= P_4_9[35];
            mult_part_out15[320] <= P_4_10[12];
            mult_part_out15[321] <= P_14_3[11];
            mult_part_out15[322] <= P_10_6[8];
            mult_part_out15[323] <= P_5_9[22];
            mult_part_out15[324] <= P_12_5[0];
            mult_part_out15[325] <= P_9_7[4];
            mult_part_out15[326] <= P_14_3[16];
            mult_part_out15[327] <= P_13_4[10];
            mult_part_out15[328] <= P_13_3[35];
            mult_part_out15[329] <= P_6_8[35];
            mult_part_out15[330] <= P_13_3[37];
            mult_part_out15[331] <= P_5_9[30];
            mult_part_out15[332] <= P_6_9[14];
            mult_part_out15[333] <= P_14_3[23];
            mult_part_out15[334] <= P_9_7[13];
            mult_part_out15[335] <= P_10_6[21];
            mult_part_out15[336] <= P_13_4[19];
            mult_part_out15[337] <= P_5_9[36];
            mult_part_out15[338] <= P_11_5[31];
            mult_part_out15[339] <= P_14_4[5];
            mult_part_out15[340] <= P_14_3[30];
            mult_part_out15[341] <= P_15_3[14];
            mult_part_out15[342] <= P_9_7[21];
            mult_part_out15[343] <= P_11_6[12];
            mult_part_out15[344] <= P_8_7[40];
            mult_part_out15[345] <= P_11_5[38];
            mult_part_out15[346] <= P_7_8[35];
            mult_part_out15[347] <= P_7_8[36];
            mult_part_out15[348] <= P_7_9[13];
            mult_part_out15[349] <= P_12_5[25];
            mult_part_out15[350] <= P_13_5[9];
            mult_part_out15[351] <= P_7_8[40];
            mult_part_out15[352] <= P_14_4[18];
            mult_part_out15[353] <= P_8_8[25];
            mult_part_out15[354] <= P_6_10[12];
            mult_part_out15[355] <= P_9_7[34];
            mult_part_out15[356] <= P_15_4[5];
            mult_part_out15[357] <= P_12_6[9];
            mult_part_out15[358] <= P_15_4[7];
            mult_part_out15[359] <= P_11_6[28];
            mult_part_out15[360] <= P_8_9[8];
            mult_part_out15[361] <= P_10_7[23];
            mult_part_out15[362] <= P_6_10[20];
            mult_part_out15[363] <= P_11_7[8];
            mult_part_out15[364] <= P_11_6[33];
            mult_part_out15[365] <= P_14_4[31];
            mult_part_out15[366] <= P_10_8[4];
            mult_part_out15[367] <= P_13_5[26];
            mult_part_out15[368] <= P_9_8[23];
            mult_part_out15[369] <= P_13_5[28];
            mult_part_out15[370] <= P_11_6[39];
            mult_part_out15[371] <= P_8_9[19];
            mult_part_out15[372] <= P_7_9[37];
            mult_part_out15[373] <= P_7_10[14];
            mult_part_out15[374] <= P_10_8[12];

            mult_part_out16[168] <= P_6_2[18];
            mult_part_out16[169] <= P_0_6[25];
            mult_part_out16[170] <= P_4_3[30];
            mult_part_out16[171] <= P_8_1[11];
            mult_part_out16[172] <= P_7_1[29];
            mult_part_out16[173] <= P_2_5[19];
            mult_part_out16[174] <= P_0_7[6];
            mult_part_out16[175] <= P_8_0[39];
            mult_part_out16[176] <= P_4_3[36];
            mult_part_out16[177] <= P_7_2[10];
            mult_part_out16[178] <= P_3_5[7];
            mult_part_out16[179] <= P_7_1[36];
            mult_part_out16[180] <= P_2_5[26];
            mult_part_out16[181] <= P_0_7[13];
            mult_part_out16[182] <= P_5_4[1];
            mult_part_out16[183] <= P_6_3[9];
            mult_part_out16[184] <= P_7_2[17];
            mult_part_out16[185] <= P_0_7[17];
            mult_part_out16[186] <= P_9_1[9];
            mult_part_out16[187] <= P_6_3[13];
            mult_part_out16[188] <= P_9_1[11];
            mult_part_out16[189] <= P_1_7[4];
            mult_part_out16[190] <= P_4_5[2];
            mult_part_out16[191] <= P_7_3[0];
            mult_part_out16[192] <= P_1_6[31];
            mult_part_out16[193] <= P_11_0[6];
            mult_part_out16[194] <= P_2_5[40];
            mult_part_out16[195] <= P_8_2[11];
            mult_part_out16[196] <= P_9_1[19];
            mult_part_out16[197] <= P_8_1[37];
            mult_part_out16[198] <= P_1_7[13];
            mult_part_out16[199] <= P_0_7[31];
            mult_part_out16[200] <= P_3_6[5];
            mult_part_out16[201] <= P_7_2[34];
            mult_part_out16[202] <= P_7_2[35];
            mult_part_out16[203] <= P_0_7[35];
            mult_part_out16[204] <= P_1_7[19];
            mult_part_out16[205] <= P_10_1[11];
            mult_part_out16[206] <= P_7_3[15];
            mult_part_out16[207] <= P_9_2[6];
            mult_part_out16[208] <= P_5_5[3];
            mult_part_out16[209] <= P_6_3[35];
            mult_part_out16[210] <= P_4_5[22];
            mult_part_out16[211] <= P_3_5[40];
            mult_part_out16[212] <= P_11_0[25];
            mult_part_out16[213] <= P_3_6[18];
            mult_part_out16[214] <= P_10_1[20];
            mult_part_out16[215] <= P_3_6[20];
            mult_part_out16[216] <= P_7_4[1];
            mult_part_out16[217] <= P_4_5[29];
            mult_part_out16[218] <= P_3_6[23];
            mult_part_out16[219] <= P_1_8[10];
            mult_part_out16[220] <= P_7_3[29];
            mult_part_out16[221] <= P_4_5[33];
            mult_part_out16[222] <= P_5_5[17];
            mult_part_out16[223] <= P_4_5[35];
            mult_part_out16[224] <= P_7_4[9];
            mult_part_out16[225] <= P_7_3[34];
            mult_part_out16[226] <= P_3_6[31];
            mult_part_out16[227] <= P_11_0[40];
            mult_part_out16[228] <= P_10_2[10];
            mult_part_out16[229] <= P_2_8[3];
            mult_part_out16[230] <= P_0_9[14];
            mult_part_out16[231] <= P_2_8[5];
            mult_part_out16[232] <= P_10_2[14];
            mult_part_out16[233] <= P_5_6[4];
            mult_part_out16[234] <= P_8_4[2];
            mult_part_out16[235] <= P_5_5[30];
            mult_part_out16[236] <= P_5_5[31];
            mult_part_out16[237] <= P_3_7[18];
            mult_part_out16[238] <= P_12_0[34];
            mult_part_out16[239] <= P_3_7[20];
            mult_part_out16[240] <= P_9_2[39];
            mult_part_out16[241] <= P_13_0[20];
            mult_part_out16[242] <= P_1_9[9];
            mult_part_out16[243] <= P_11_1[32];
            mult_part_out16[244] <= P_7_5[5];
            mult_part_out16[245] <= P_4_6[33];
            mult_part_out16[246] <= P_11_2[11];
            mult_part_out16[247] <= P_7_4[32];
            mult_part_out16[248] <= P_12_1[20];
            mult_part_out16[249] <= P_3_7[30];
            mult_part_out16[250] <= P_7_5[11];
            mult_part_out16[251] <= P_9_3[26];
            mult_part_out16[252] <= P_14_0[14];
            mult_part_out16[253] <= P_10_3[11];
            mult_part_out16[254] <= P_0_10[14];
            mult_part_out16[255] <= P_10_3[13];
            mult_part_out16[256] <= P_8_5[0];
            mult_part_out16[257] <= P_14_0[19];
            mult_part_out16[258] <= P_13_1[13];
            mult_part_out16[259] <= P_6_6[13];
            mult_part_out16[260] <= P_12_2[8];
            mult_part_out16[261] <= P_13_1[16];
            mult_part_out16[262] <= P_3_8[19];
            mult_part_out16[263] <= P_6_6[17];
            mult_part_out16[264] <= P_8_4[32];
            mult_part_out16[265] <= P_5_6[36];
            mult_part_out16[266] <= P_15_0[11];
            mult_part_out16[267] <= P_8_5[11];
            mult_part_out16[268] <= P_4_8[8];
            mult_part_out16[269] <= P_13_1[24];
            mult_part_out16[270] <= P_14_1[8];
            mult_part_out16[271] <= P_14_0[33];
            mult_part_out16[272] <= P_1_10[15];
            mult_part_out16[273] <= P_10_3[31];
            mult_part_out16[274] <= P_2_9[24];
            mult_part_out16[275] <= P_6_6[29];
            mult_part_out16[276] <= P_4_7[40];
            mult_part_out16[277] <= P_6_7[7];
            mult_part_out16[278] <= P_2_9[28];
            mult_part_out16[279] <= P_6_7[9];
            mult_part_out16[280] <= P_9_4[31];
            mult_part_out16[281] <= P_13_1[36];
            mult_part_out16[282] <= P_14_1[20];
            mult_part_out16[283] <= P_2_9[33];
            mult_part_out16[284] <= P_8_5[28];
            mult_part_out16[285] <= P_9_4[36];
            mult_part_out16[286] <= P_2_9[36];
            mult_part_out16[287] <= P_5_7[34];
            mult_part_out16[288] <= P_12_3[12];
            mult_part_out16[289] <= P_14_2[3];
            mult_part_out16[290] <= P_2_10[16];
            mult_part_out16[291] <= P_11_3[32];
            mult_part_out16[292] <= P_3_10[1];
            mult_part_out16[293] <= P_5_8[16];
            mult_part_out16[294] <= P_7_7[7];
            mult_part_out16[295] <= P_11_3[36];
            mult_part_out16[296] <= P_9_5[23];
            mult_part_out16[297] <= P_6_8[3];
            mult_part_out16[298] <= P_10_4[32];
            mult_part_out16[299] <= P_5_8[22];
            mult_part_out16[300] <= P_13_3[7];
            mult_part_out16[301] <= P_12_4[1];
            mult_part_out16[302] <= P_10_5[12];
            mult_part_out16[303] <= P_4_9[19];
            mult_part_out16[304] <= P_9_5[31];
            mult_part_out16[305] <= P_13_3[12];
            mult_part_out16[306] <= P_13_2[37];
            mult_part_out16[307] <= P_11_5[0];
            mult_part_out16[308] <= P_10_5[18];
            mult_part_out16[309] <= P_9_5[36];
            mult_part_out16[310] <= P_13_3[17];
            mult_part_out16[311] <= P_5_9[10];
            mult_part_out16[312] <= P_11_4[29];
            mult_part_out16[313] <= P_4_9[29];
            mult_part_out16[314] <= P_10_5[24];
            mult_part_out16[315] <= P_4_9[31];
            mult_part_out16[316] <= P_14_2[30];
            mult_part_out16[317] <= P_7_8[6];
            mult_part_out16[318] <= P_14_3[8];
            mult_part_out16[319] <= P_14_3[9];
            mult_part_out16[320] <= P_5_9[19];
            mult_part_out16[321] <= P_6_8[27];
            mult_part_out16[322] <= P_14_3[12];
            mult_part_out16[323] <= P_11_4[40];
            mult_part_out16[324] <= P_10_5[34];
            mult_part_out16[325] <= P_8_7[21];
            mult_part_out16[326] <= P_9_7[5];
            mult_part_out16[327] <= P_15_3[0];
            mult_part_out16[328] <= P_5_9[27];
            mult_part_out16[329] <= P_5_9[28];
            mult_part_out16[330] <= P_10_5[40];
            mult_part_out16[331] <= P_11_6[0];
            mult_part_out16[332] <= P_14_3[22];
            mult_part_out16[333] <= P_8_7[29];
            mult_part_out16[334] <= P_9_6[37];
            mult_part_out16[335] <= P_13_4[18];
            mult_part_out16[336] <= P_11_5[29];
            mult_part_out16[337] <= P_9_7[16];
            mult_part_out16[338] <= P_10_7[0];
            mult_part_out16[339] <= P_11_5[32];
            mult_part_out16[340] <= P_11_6[9];
            mult_part_out16[341] <= P_5_9[40];
            mult_part_out16[342] <= P_7_9[7];
            mult_part_out16[343] <= P_13_5[2];
            mult_part_out16[344] <= P_6_10[2];
            mult_part_out16[345] <= P_10_6[31];
            mult_part_out16[346] <= P_5_10[21];
            mult_part_out16[347] <= P_10_7[9];
            mult_part_out16[348] <= P_10_6[34];
            mult_part_out16[349] <= P_14_3[39];
            mult_part_out16[350] <= P_6_9[32];
            mult_part_out16[351] <= P_13_4[34];
            mult_part_out16[352] <= P_10_7[14];
            mult_part_out16[353] <= P_10_6[39];
            mult_part_out16[354] <= P_13_5[13];
            mult_part_out16[355] <= P_7_9[20];
            mult_part_out16[356] <= P_12_6[8];
            mult_part_out16[357] <= P_9_8[12];

            mult_part_out17[170] <= P_7_1[27];
            mult_part_out17[171] <= P_0_6[27];
            mult_part_out17[172] <= P_9_0[19];
            mult_part_out17[173] <= P_1_6[12];
            mult_part_out17[174] <= P_2_5[20];
            mult_part_out17[175] <= P_8_1[15];
            mult_part_out17[176] <= P_7_2[9];
            mult_part_out17[177] <= P_1_5[40];
            mult_part_out17[178] <= P_9_1[1];
            mult_part_out17[179] <= P_10_0[9];
            mult_part_out17[180] <= P_9_0[27];
            mult_part_out17[181] <= P_8_1[21];
            mult_part_out17[182] <= P_9_0[29];
            mult_part_out17[183] <= P_5_3[26];
            mult_part_out17[184] <= P_3_4[37];
            mult_part_out17[185] <= P_9_0[32];
            mult_part_out17[186] <= P_9_0[33];
            mult_part_out17[187] <= P_0_7[19];
            mult_part_out17[188] <= P_7_2[21];
            mult_part_out17[189] <= P_7_2[22];
            mult_part_out17[190] <= P_5_3[33];
            mult_part_out17[191] <= P_2_5[37];
            mult_part_out17[192] <= P_4_5[4];
            mult_part_out17[193] <= P_0_8[1];
            mult_part_out17[194] <= P_4_4[30];
            mult_part_out17[195] <= P_0_8[3];
            mult_part_out17[196] <= P_1_6[35];
            mult_part_out17[197] <= P_10_1[3];
            mult_part_out17[198] <= P_4_5[10];
            mult_part_out17[199] <= P_3_6[4];
            mult_part_out17[200] <= P_4_5[12];
            mult_part_out17[201] <= P_8_2[17];
            mult_part_out17[202] <= P_3_6[7];
            mult_part_out17[203] <= P_4_5[15];
            mult_part_out17[204] <= P_12_0[0];
            mult_part_out17[205] <= P_2_7[3];
            mult_part_out17[206] <= P_7_2[39];
            mult_part_out17[207] <= P_9_1[30];
            mult_part_out17[208] <= P_10_1[14];
            mult_part_out17[209] <= P_8_2[25];
            mult_part_out17[210] <= P_9_2[9];
            mult_part_out17[211] <= P_11_0[24];
            mult_part_out17[212] <= P_7_3[21];
            mult_part_out17[213] <= P_1_7[28];
            mult_part_out17[214] <= P_11_1[3];
            mult_part_out17[215] <= P_4_5[27];
            mult_part_out17[216] <= P_8_2[32];
            mult_part_out17[217] <= P_9_1[40];
            mult_part_out17[218] <= P_5_5[13];
            mult_part_out17[219] <= P_5_5[14];
            mult_part_out17[220] <= P_8_3[12];
            mult_part_out17[221] <= P_4_6[9];
            mult_part_out17[222] <= P_2_7[20];
            mult_part_out17[223] <= P_11_0[36];
            mult_part_out17[224] <= P_8_2[40];
            mult_part_out17[225] <= P_10_2[7];
            mult_part_out17[226] <= P_9_3[1];
            mult_part_out17[227] <= P_11_1[16];
            mult_part_out17[228] <= P_7_4[13];
            mult_part_out17[229] <= P_5_6[0];
            mult_part_out17[230] <= P_4_6[18];
            mult_part_out17[231] <= P_13_0[10];
            mult_part_out17[232] <= P_2_8[6];
            mult_part_out17[233] <= P_2_8[7];
            mult_part_out17[234] <= P_2_7[32];
            mult_part_out17[235] <= P_2_7[33];
            mult_part_out17[236] <= P_11_1[25];
            mult_part_out17[237] <= P_7_4[22];
            mult_part_out17[238] <= P_14_0[0];
            mult_part_out17[239] <= P_5_6[10];
            mult_part_out17[240] <= P_4_7[4];
            mult_part_out17[241] <= P_12_0[37];
            mult_part_out17[242] <= P_2_7[40];
            mult_part_out17[243] <= P_7_4[28];
            mult_part_out17[244] <= P_5_6[15];
            mult_part_out17[245] <= P_11_1[34];
            mult_part_out17[246] <= P_9_3[21];
            mult_part_out17[247] <= P_1_9[14];
            mult_part_out17[248] <= P_3_8[5];
            mult_part_out17[249] <= P_5_6[20];
            mult_part_out17[250] <= P_1_9[17];
            mult_part_out17[251] <= P_1_9[18];
            mult_part_out17[252] <= P_2_9[2];
            mult_part_out17[253] <= P_5_7[0];
            mult_part_out17[254] <= P_5_6[25];
            mult_part_out17[255] <= P_8_4[23];
            mult_part_out17[256] <= P_5_7[3];
            mult_part_out17[257] <= P_6_6[11];
            mult_part_out17[258] <= P_2_9[8];
            mult_part_out17[259] <= P_13_1[14];
            mult_part_out17[260] <= P_2_9[10];
            mult_part_out17[261] <= P_5_6[32];
            mult_part_out17[262] <= P_6_5[40];
            mult_part_out17[263] <= P_8_4[31];
            mult_part_out17[264] <= P_15_0[9];
            mult_part_out17[265] <= P_14_0[27];
            mult_part_out17[266] <= P_2_8[40];
            mult_part_out17[267] <= P_14_1[5];
            mult_part_out17[268] <= P_3_9[1];
            mult_part_out17[269] <= P_4_8[9];
            mult_part_out17[270] <= P_15_0[15];
            mult_part_out17[271] <= P_3_9[4];
            mult_part_out17[272] <= P_11_2[37];
            mult_part_out17[273] <= P_8_5[17];
            mult_part_out17[274] <= P_3_8[31];
            mult_part_out17[275] <= P_10_4[9];
            mult_part_out17[276] <= P_9_4[27];
            mult_part_out17[277] <= P_3_9[10];
            mult_part_out17[278] <= P_13_2[9];
            mult_part_out17[279] <= P_15_0[24];
            mult_part_out17[280] <= P_15_1[1];
            mult_part_out17[281] <= P_2_9[31];
            mult_part_out17[282] <= P_2_10[8];
            mult_part_out17[283] <= P_6_7[13];
            mult_part_out17[284] <= P_13_1[39];
            mult_part_out17[285] <= P_6_6[39];
            mult_part_out17[286] <= P_8_5[30];
            mult_part_out17[287] <= P_8_5[31];
            mult_part_out17[288] <= P_3_9[21];
            mult_part_out17[289] <= P_10_4[23];
            mult_part_out17[290] <= P_12_3[14];
            mult_part_out17[291] <= P_8_6[11];
            mult_part_out17[292] <= P_12_3[16];
            mult_part_out17[293] <= P_7_7[6];
            mult_part_out17[294] <= P_4_9[10];
            mult_part_out17[295] <= P_13_3[2];
            mult_part_out17[296] <= P_2_10[22];
            mult_part_out17[297] <= P_12_3[21];
            mult_part_out17[298] <= P_6_8[4];
            mult_part_out17[299] <= P_6_7[29];
            mult_part_out17[300] <= P_7_6[37];
            mult_part_out17[301] <= P_9_6[4];
            mult_part_out17[302] <= P_5_8[25];
            mult_part_out17[303] <= P_12_4[3];
            mult_part_out17[304] <= P_3_10[13];
            mult_part_out17[305] <= P_12_3[29];
            mult_part_out17[306] <= P_7_7[19];
            mult_part_out17[307] <= P_8_7[3];
            mult_part_out17[308] <= P_3_10[17];
            mult_part_out17[309] <= P_14_2[23];
            mult_part_out17[310] <= P_9_6[13];
            mult_part_out17[311] <= P_9_5[38];
            mult_part_out17[312] <= P_7_7[25];
            mult_part_out17[313] <= P_14_3[3];
            mult_part_out17[314] <= P_10_6[0];
            mult_part_out17[315] <= P_8_6[35];
            mult_part_out17[316] <= P_4_9[32];
            mult_part_out17[317] <= P_13_3[24];
            mult_part_out17[318] <= P_11_4[35];
            mult_part_out17[319] <= P_15_2[16];
            mult_part_out17[320] <= P_15_2[17];
            mult_part_out17[321] <= P_10_6[7];
            mult_part_out17[322] <= P_15_2[19];
            mult_part_out17[323] <= P_13_3[30];
            mult_part_out17[324] <= P_8_7[20];
            mult_part_out17[325] <= P_13_4[8];
            mult_part_out17[326] <= P_9_6[29];
            mult_part_out17[327] <= P_15_2[24];
            mult_part_out17[328] <= P_12_4[28];
            mult_part_out17[329] <= P_6_9[11];
            mult_part_out17[330] <= P_14_3[20];
            mult_part_out17[331] <= P_8_7[27];
            mult_part_out17[332] <= P_8_7[28];
            mult_part_out17[333] <= P_6_8[39];
            mult_part_out17[334] <= P_5_10[9];
            mult_part_out17[335] <= P_12_5[11];
            mult_part_out17[336] <= P_6_9[18];
            mult_part_out17[337] <= P_14_3[27];
            mult_part_out17[338] <= P_10_6[24];
            mult_part_out17[339] <= P_15_3[12];
            mult_part_out17[340] <= P_9_7[19];
            mult_part_out17[341] <= P_11_6[10];
            mult_part_out17[342] <= P_12_5[18];
            mult_part_out17[343] <= P_9_7[22];
            mult_part_out17[344] <= P_5_10[19];
            mult_part_out17[345] <= P_11_6[14];
            mult_part_out17[346] <= P_13_4[29];
            mult_part_out17[347] <= P_6_9[29];
            mult_part_out17[348] <= P_6_9[30];
            mult_part_out17[349] <= P_15_3[22];
            mult_part_out17[350] <= P_7_9[15];
            mult_part_out17[351] <= P_14_4[17];

            mult_part_out18[187] <= P_11_0[0];
            mult_part_out18[188] <= P_3_5[17];
            mult_part_out18[189] <= P_2_5[35];
            mult_part_out18[190] <= P_5_4[9];
            mult_part_out18[191] <= P_1_7[6];
            mult_part_out18[192] <= P_0_8[0];
            mult_part_out18[193] <= P_8_1[33];
            mult_part_out18[194] <= P_0_8[2];
            mult_part_out18[195] <= P_11_0[8];
            mult_part_out18[196] <= P_7_2[29];
            mult_part_out18[197] <= P_7_2[30];
            mult_part_out18[198] <= P_6_4[0];
            mult_part_out18[199] <= P_8_1[39];
            mult_part_out18[200] <= P_8_2[16];
            mult_part_out18[201] <= P_4_5[13];
            mult_part_out18[202] <= P_5_4[21];
            mult_part_out18[203] <= P_11_0[16];
            mult_part_out18[204] <= P_6_3[30];
            mult_part_out18[205] <= P_3_6[10];
            mult_part_out18[206] <= P_10_1[12];
            mult_part_out18[207] <= P_7_3[16];
            mult_part_out18[208] <= P_6_3[34];
            mult_part_out18[209] <= P_3_6[14];
            mult_part_out18[210] <= P_5_5[5];
            mult_part_out18[211] <= P_11_1[0];
            mult_part_out18[212] <= P_11_1[1];
            mult_part_out18[213] <= P_9_2[12];
            mult_part_out18[214] <= P_11_0[27];
            mult_part_out18[215] <= P_2_6[37];
            mult_part_out18[216] <= P_6_4[18];
            mult_part_out18[217] <= P_1_7[32];
            mult_part_out18[218] <= P_6_4[20];
            mult_part_out18[219] <= P_5_4[38];
            mult_part_out18[220] <= P_10_2[2];
            mult_part_out18[221] <= P_6_4[23];
            mult_part_out18[222] <= P_0_8[30];
            mult_part_out18[223] <= P_5_5[18];
            mult_part_out18[224] <= P_3_7[5];
            mult_part_out18[225] <= P_3_7[6];
            mult_part_out18[226] <= P_1_8[17];
            mult_part_out18[227] <= P_7_4[12];
            mult_part_out18[228] <= P_6_5[6];
            mult_part_out18[229] <= P_1_8[20];
            mult_part_out18[230] <= P_5_5[25];
            mult_part_out18[231] <= P_5_5[26];
            mult_part_out18[232] <= P_4_6[20];
            mult_part_out18[233] <= P_2_7[31];
            mult_part_out18[234] <= P_11_1[23];
            mult_part_out18[235] <= P_0_9[19];
            mult_part_out18[236] <= P_12_0[32];
            mult_part_out18[237] <= P_5_5[32];
            mult_part_out18[238] <= P_1_8[29];
            mult_part_out18[239] <= P_7_4[24];
            mult_part_out18[240] <= P_0_10[0];
            mult_part_out18[241] <= P_4_7[5];
            mult_part_out18[242] <= P_6_5[20];
            mult_part_out18[243] <= P_4_7[7];
            mult_part_out18[244] <= P_12_1[16];
            mult_part_out18[245] <= P_5_6[16];
            mult_part_out18[246] <= P_10_2[28];
            mult_part_out18[247] <= P_6_6[1];
            mult_part_out18[248] <= P_13_1[3];
            mult_part_out18[249] <= P_10_2[31];
            mult_part_out18[250] <= P_9_3[25];
            mult_part_out18[251] <= P_6_6[5];
            mult_part_out18[252] <= P_0_10[12];
            mult_part_out18[253] <= P_0_9[37];
            mult_part_out18[254] <= P_7_4[39];
            mult_part_out18[255] <= P_9_4[6];
            mult_part_out18[256] <= P_2_9[6];
            mult_part_out18[257] <= P_7_5[18];
            mult_part_out18[258] <= P_11_2[23];
            mult_part_out18[259] <= P_2_9[9];
            mult_part_out18[260] <= P_12_1[32];
            mult_part_out18[261] <= P_11_3[2];
            mult_part_out18[262] <= P_1_10[5];
            mult_part_out18[263] <= P_10_3[21];
            mult_part_out18[264] <= P_7_6[1];
            mult_part_out18[265] <= P_14_1[3];
            mult_part_out18[266] <= P_10_3[24];
            mult_part_out18[267] <= P_1_10[10];
            mult_part_out18[268] <= P_7_5[29];
            mult_part_out18[269] <= P_9_4[20];
            mult_part_out18[270] <= P_9_4[21];
            mult_part_out18[271] <= P_4_8[11];
            mult_part_out18[272] <= P_12_2[20];
            mult_part_out18[273] <= P_4_8[13];
            mult_part_out18[274] <= P_7_5[35];
            mult_part_out18[275] <= P_13_2[6];
            mult_part_out18[276] <= P_13_2[7];
            mult_part_out18[277] <= P_9_4[28];
            mult_part_out18[278] <= P_14_1[16];
            mult_part_out18[279] <= P_2_9[29];
            mult_part_out18[280] <= P_2_10[6];
            mult_part_out18[281] <= P_13_2[12];
            mult_part_out18[282] <= P_10_3[40];
            mult_part_out18[283] <= P_11_3[24];
            mult_part_out18[284] <= P_6_7[14];
            mult_part_out18[285] <= P_8_6[5];
            mult_part_out18[286] <= P_5_7[33];
            mult_part_out18[287] <= P_7_6[24];
            mult_part_out18[288] <= P_11_3[29];
            mult_part_out18[289] <= P_7_7[2];
            mult_part_out18[290] <= P_3_9[23];
            mult_part_out18[291] <= P_2_10[17];
            mult_part_out18[292] <= P_13_2[23];
            mult_part_out18[293] <= P_13_3[0];
            mult_part_out18[294] <= P_13_2[25];
            mult_part_out18[295] <= P_8_6[15];
            mult_part_out18[296] <= P_4_9[12];
            mult_part_out18[297] <= P_4_8[37];
            mult_part_out18[298] <= P_5_8[21];
            mult_part_out18[299] <= P_4_8[39];
            mult_part_out18[300] <= P_8_6[20];
            mult_part_out18[301] <= P_10_5[11];
            mult_part_out18[302] <= P_11_4[19];
            mult_part_out18[303] <= P_8_6[23];
            mult_part_out18[304] <= P_10_4[38];
            mult_part_out18[305] <= P_6_8[11];
            mult_part_out18[306] <= P_13_3[13];
            mult_part_out18[307] <= P_12_3[31];
            mult_part_out18[308] <= P_5_9[7];
            mult_part_out18[309] <= P_8_6[29];
            mult_part_out18[310] <= P_5_8[33];
            mult_part_out18[311] <= P_8_6[31];
            mult_part_out18[312] <= P_6_8[18];
            mult_part_out18[313] <= P_10_5[23];
            mult_part_out18[314] <= P_11_4[31];
            mult_part_out18[315] <= P_10_6[1];
            mult_part_out18[316] <= P_11_5[9];
            mult_part_out18[317] <= P_13_4[0];
            mult_part_out18[318] <= P_6_9[0];
            mult_part_out18[319] <= P_10_6[5];
            mult_part_out18[320] <= P_7_8[9];
            mult_part_out18[321] <= P_10_5[31];
            mult_part_out18[322] <= P_6_8[28];
            mult_part_out18[323] <= P_8_7[19];
            mult_part_out18[324] <= P_10_6[10];
            mult_part_out18[325] <= P_10_5[35];
            mult_part_out18[326] <= P_10_6[12];
            mult_part_out18[327] <= P_14_3[17];
            mult_part_out18[328] <= P_11_5[21];
            mult_part_out18[329] <= P_8_8[1];
            mult_part_out18[330] <= P_6_8[36];
            mult_part_out18[331] <= P_12_4[31];
            mult_part_out18[332] <= P_11_6[1];
            mult_part_out18[333] <= P_9_6[36];
            mult_part_out18[334] <= P_14_3[24];
            mult_part_out18[335] <= P_15_3[8];
            mult_part_out18[336] <= P_5_10[11];
            mult_part_out18[337] <= P_8_8[9];
            mult_part_out18[338] <= P_14_3[28];
            mult_part_out18[339] <= P_11_6[8];
            mult_part_out18[340] <= P_7_9[5];

            mult_part_out19[192] <= P_9_1[15];
            mult_part_out19[193] <= P_4_5[5];
            mult_part_out19[194] <= P_11_0[7];
            mult_part_out19[195] <= P_8_1[35];
            mult_part_out19[196] <= P_7_3[5];
            mult_part_out19[197] <= P_3_6[2];
            mult_part_out19[198] <= P_6_3[24];
            mult_part_out19[199] <= P_4_4[35];
            mult_part_out19[200] <= P_9_1[23];
            mult_part_out19[201] <= P_1_6[40];
            mult_part_out19[202] <= P_6_3[28];
            mult_part_out19[203] <= P_4_4[39];
            mult_part_out19[204] <= P_10_1[10];
            mult_part_out19[205] <= P_9_2[4];
            mult_part_out19[206] <= P_6_4[8];
            mult_part_out19[207] <= P_0_8[15];
            mult_part_out19[208] <= P_8_2[24];
            mult_part_out19[209] <= P_10_0[39];
            mult_part_out19[210] <= P_8_2[26];
            mult_part_out19[211] <= P_12_0[7];
            mult_part_out19[212] <= P_8_3[4];
            mult_part_out19[213] <= P_2_7[11];
            mult_part_out19[214] <= P_7_3[23];
            mult_part_out19[215] <= P_0_8[23];
            mult_part_out19[216] <= P_1_7[31];
            mult_part_out19[217] <= P_8_2[33];
            mult_part_out19[218] <= P_10_1[24];
            mult_part_out19[219] <= P_3_6[24];
            mult_part_out19[220] <= P_5_5[15];
            mult_part_out19[221] <= P_3_7[2];
            mult_part_out19[222] <= P_8_2[38];
            mult_part_out19[223] <= P_3_6[28];
            mult_part_out19[224] <= P_6_5[2];
            mult_part_out19[225] <= P_3_6[30];
            mult_part_out19[226] <= P_4_5[38];
            mult_part_out19[227] <= P_3_6[32];
            mult_part_out19[228] <= P_1_8[19];
            mult_part_out19[229] <= P_2_7[27];
            mult_part_out19[230] <= P_0_8[38];
            mult_part_out19[231] <= P_5_6[2];
            mult_part_out19[232] <= P_5_6[3];
            mult_part_out19[233] <= P_9_2[32];
            mult_part_out19[234] <= P_5_6[5];
            mult_part_out19[235] <= P_10_2[17];
            mult_part_out19[236] <= P_6_4[38];
            mult_part_out19[237] <= P_9_3[12];
            mult_part_out19[238] <= P_9_2[37];
            mult_part_out19[239] <= P_13_0[18];
            mult_part_out19[240] <= P_4_6[28];
            mult_part_out19[241] <= P_5_5[36];
            mult_part_out19[242] <= P_5_6[13];
            mult_part_out19[243] <= P_6_5[21];
            mult_part_out19[244] <= P_11_2[9];
            mult_part_out19[245] <= P_10_2[27];
            mult_part_out19[246] <= P_8_3[38];
            mult_part_out19[247] <= P_10_3[5];
            mult_part_out19[248] <= P_7_4[33];
            mult_part_out19[249] <= P_1_9[16];
            mult_part_out19[250] <= P_2_8[24];
            mult_part_out19[251] <= P_14_0[13];
            mult_part_out19[252] <= P_3_7[33];
            mult_part_out19[253] <= P_9_3[28];
            mult_part_out19[254] <= P_13_0[33];
            mult_part_out19[255] <= P_5_7[2];
            mult_part_out19[256] <= P_11_2[21];
            mult_part_out19[257] <= P_12_2[5];
            mult_part_out19[258] <= P_6_5[36];
            mult_part_out19[259] <= P_3_7[40];
            mult_part_out19[260] <= P_4_8[0];
            mult_part_out19[261] <= P_8_4[29];
            mult_part_out19[262] <= P_8_4[30];
            mult_part_out19[263] <= P_12_2[11];
            mult_part_out19[264] <= P_13_1[19];
            mult_part_out19[265] <= P_2_8[39];
            mult_part_out19[266] <= P_0_10[26];
            mult_part_out19[267] <= P_6_6[21];
            mult_part_out19[268] <= P_3_8[25];
            mult_part_out19[269] <= P_15_0[14];
            mult_part_out19[270] <= P_3_9[3];
            mult_part_out19[271] <= P_14_1[9];
            mult_part_out19[272] <= P_13_1[27];
            mult_part_out19[273] <= P_5_7[20];
            mult_part_out19[274] <= P_9_4[25];
            mult_part_out19[275] <= P_7_6[12];
            mult_part_out19[276] <= P_15_0[21];
            mult_part_out19[277] <= P_15_0[22];
            mult_part_out19[278] <= P_7_5[39];
            mult_part_out19[279] <= P_10_3[37];
            mult_part_out19[280] <= P_7_6[17];
            mult_part_out19[281] <= P_6_7[11];
            mult_part_out19[282] <= P_12_2[30];
            mult_part_out19[283] <= P_8_6[3];
            mult_part_out19[284] <= P_3_9[17];
            mult_part_out19[285] <= P_8_5[29];
            mult_part_out19[286] <= P_4_9[2];
            mult_part_out19[287] <= P_9_4[38];
            mult_part_out19[288] <= P_9_4[39];
            mult_part_out19[289] <= P_14_1[27];
            mult_part_out19[290] <= P_12_2[38];
            mult_part_out19[291] <= P_5_7[38];
            mult_part_out19[292] <= P_8_5[36];
            mult_part_out19[293] <= P_4_8[33];
            mult_part_out19[294] <= P_15_1[15];
            mult_part_out19[295] <= P_12_3[19];
            mult_part_out19[296] <= P_10_4[30];
            mult_part_out19[297] <= P_14_2[11];
            mult_part_out19[298] <= P_12_3[22];
            mult_part_out19[299] <= P_10_5[9];
            mult_part_out19[300] <= P_12_4[0];
            mult_part_out19[301] <= P_5_8[24];
            mult_part_out19[302] <= P_13_3[9];
            mult_part_out19[303] <= P_13_2[34];
            mult_part_out19[304] <= P_7_7[17];
            mult_part_out19[305] <= P_9_5[32];
            mult_part_out19[306] <= P_2_10[32];
            mult_part_out19[307] <= P_10_5[17];
            mult_part_out19[308] <= P_8_6[28];
            mult_part_out19[309] <= P_9_6[12];
            mult_part_out19[310] <= P_8_6[30];
            mult_part_out19[311] <= P_9_6[14];
            mult_part_out19[312] <= P_7_8[1];
            mult_part_out19[313] <= P_8_7[9];
            mult_part_out19[314] <= P_4_10[6];
            mult_part_out19[315] <= P_14_3[5];
            mult_part_out19[316] <= P_11_4[33];
            mult_part_out19[317] <= P_14_2[31];
            mult_part_out19[318] <= P_3_10[27];
            mult_part_out19[319] <= P_6_9[1];
            mult_part_out19[320] <= P_12_4[20];
            mult_part_out19[321] <= P_14_2[35];
            mult_part_out19[322] <= P_13_4[5];
            mult_part_out19[323] <= P_11_5[16];
            mult_part_out19[324] <= P_6_9[6];
            mult_part_out19[325] <= P_12_5[1];
            mult_part_out19[326] <= P_15_2[23];
            mult_part_out19[327] <= P_6_9[9];

            mult_part_out20[204] <= P_8_2[20];
            mult_part_out20[205] <= P_9_1[28];
            mult_part_out20[206] <= P_5_5[1];
            mult_part_out20[207] <= P_2_6[29];
            mult_part_out20[208] <= P_0_7[40];
            mult_part_out20[209] <= P_9_2[8];
            mult_part_out20[210] <= P_1_8[1];
            mult_part_out20[211] <= P_4_5[23];
            mult_part_out20[212] <= P_10_1[18];
            mult_part_out20[213] <= P_2_6[35];
            mult_part_out20[214] <= P_8_3[6];
            mult_part_out20[215] <= P_9_2[14];
            mult_part_out20[216] <= P_1_8[7];
            mult_part_out20[217] <= P_3_6[22];
            mult_part_out20[218] <= P_4_6[6];
            mult_part_out20[219] <= P_0_9[3];
            mult_part_out20[220] <= P_7_4[5];
            mult_part_out20[221] <= P_7_4[6];
            mult_part_out20[222] <= P_13_0[1];
            mult_part_out20[223] <= P_11_1[12];
            mult_part_out20[224] <= P_4_6[12];
            mult_part_out20[225] <= P_4_6[13];
            mult_part_out20[226] <= P_7_3[35];
            mult_part_out20[227] <= P_4_5[39];
            mult_part_out20[228] <= P_10_1[34];
            mult_part_out20[229] <= P_7_3[38];
            mult_part_out20[230] <= P_6_4[32];
            mult_part_out20[231] <= P_10_2[13];
            mult_part_out20[232] <= P_9_2[31];
            mult_part_out20[233] <= P_5_5[28];
            mult_part_out20[234] <= P_4_6[22];
            mult_part_out20[235] <= P_12_1[7];
            mult_part_out20[236] <= P_2_7[34];
            mult_part_out20[237] <= P_6_4[39];
            mult_part_out20[238] <= P_9_3[13];
            mult_part_out20[239] <= P_12_1[11];
            mult_part_out20[240] <= P_11_1[29];
            mult_part_out20[241] <= P_4_6[29];
            mult_part_out20[242] <= P_11_1[31];
            mult_part_out20[243] <= P_3_7[24];
            mult_part_out20[244] <= P_8_3[36];
            mult_part_out20[245] <= P_1_9[12];
            mult_part_out20[246] <= P_8_4[14];
            mult_part_out20[247] <= P_8_4[15];
            mult_part_out20[248] <= P_5_6[19];
            mult_part_out20[249] <= P_6_5[27];
            mult_part_out20[250] <= P_0_9[34];
            mult_part_out20[251] <= P_0_10[11];
            mult_part_out20[252] <= P_4_6[40];
            mult_part_out20[253] <= P_7_5[14];
            mult_part_out20[254] <= P_13_1[9];
            mult_part_out20[255] <= P_7_5[16];
            mult_part_out20[256] <= P_0_9[40];
            mult_part_out20[257] <= P_3_8[14];
            mult_part_out20[258] <= P_8_5[2];
            mult_part_out20[259] <= P_14_0[21];
            mult_part_out20[260] <= P_8_4[28];
            mult_part_out20[261] <= P_4_7[25];
            mult_part_out20[262] <= P_1_9[29];
            mult_part_out20[263] <= P_13_1[18];
            mult_part_out20[264] <= P_9_4[15];
            mult_part_out20[265] <= P_12_2[13];
            mult_part_out20[266] <= P_8_4[34];
            mult_part_out20[267] <= P_10_4[1];
            mult_part_out20[268] <= P_14_1[6];
            mult_part_out20[269] <= P_14_1[7];
            mult_part_out20[270] <= P_6_6[24];
            mult_part_out20[271] <= P_0_10[31];
            mult_part_out20[272] <= P_7_5[33];
            mult_part_out20[273] <= P_1_9[40];
            mult_part_out20[274] <= P_2_10[0];
            mult_part_out20[275] <= P_6_7[5];
            mult_part_out20[276] <= P_13_1[31];
            mult_part_out20[277] <= P_12_3[1];
            mult_part_out20[278] <= P_3_8[35];
            mult_part_out20[279] <= P_15_1[0];
            mult_part_out20[280] <= P_12_2[28];
            mult_part_out20[281] <= P_15_1[2];
            mult_part_out20[282] <= P_12_3[6];
            mult_part_out20[283] <= P_9_5[10];
            mult_part_out20[284] <= P_2_9[34];
            mult_part_out20[285] <= P_4_8[25];
            mult_part_out20[286] <= P_4_8[26];
            mult_part_out20[287] <= P_11_3[28];
            mult_part_out20[288] <= P_9_5[15];
            mult_part_out20[289] <= P_11_4[6];
            mult_part_out20[290] <= P_6_7[20];
            mult_part_out20[291] <= P_13_2[22];
            mult_part_out20[292] <= P_11_4[9];
            mult_part_out20[293] <= P_3_9[26];
            mult_part_out20[294] <= P_14_2[8];
            mult_part_out20[295] <= P_11_4[12];
            mult_part_out20[296] <= P_7_7[9];
            mult_part_out20[297] <= P_3_10[6];
            mult_part_out20[298] <= P_7_7[11];
            mult_part_out20[299] <= P_13_2[30];
            mult_part_out20[300] <= P_7_7[13];
            mult_part_out20[301] <= P_6_7[31];
            mult_part_out20[302] <= P_10_4[36];
            mult_part_out20[303] <= P_6_7[33];
            mult_part_out20[304] <= P_2_10[30];
            mult_part_out20[305] <= P_14_2[19];
            mult_part_out20[306] <= P_11_4[23];
            mult_part_out20[307] <= P_9_5[34];
            mult_part_out20[308] <= P_9_6[11];
            mult_part_out20[309] <= P_6_8[15];
            mult_part_out20[310] <= P_3_10[19];
            mult_part_out20[311] <= P_7_7[24];
            mult_part_out20[312] <= P_13_3[19];
            mult_part_out20[313] <= P_8_6[33];
            mult_part_out20[314] <= P_14_2[28];
            mult_part_out20[315] <= P_5_9[14];
            mult_part_out20[316] <= P_8_7[12];
            mult_part_out20[317] <= P_11_4[34];
            mult_part_out20[318] <= P_11_5[11];
            mult_part_out20[319] <= P_14_2[33];
            mult_part_out20[320] <= P_14_3[10];
            mult_part_out20[321] <= P_13_4[4];
            mult_part_out20[322] <= P_12_4[22];
            mult_part_out20[323] <= P_6_9[5];

            mult_part_out21[216] <= P_11_1[5];
            mult_part_out21[217] <= P_5_5[12];
            mult_part_out21[218] <= P_1_7[33];
            mult_part_out21[219] <= P_1_7[34];
            mult_part_out21[220] <= P_12_0[16];
            mult_part_out21[221] <= P_5_4[40];
            mult_part_out21[222] <= P_1_8[13];
            mult_part_out21[223] <= P_12_0[19];
            mult_part_out21[224] <= P_5_5[19];
            mult_part_out21[225] <= P_12_0[21];
            mult_part_out21[226] <= P_3_7[7];
            mult_part_out21[227] <= P_12_0[23];
            mult_part_out21[228] <= P_12_0[24];
            mult_part_out21[229] <= P_0_9[13];
            mult_part_out21[230] <= P_7_4[15];
            mult_part_out21[231] <= P_6_5[9];
            mult_part_out21[232] <= P_5_5[27];
            mult_part_out21[233] <= P_11_1[22];
            mult_part_out21[234] <= P_7_4[19];
            mult_part_out21[235] <= P_4_6[23];
            mult_part_out21[236] <= P_0_9[20];
            mult_part_out21[237] <= P_4_6[25];
            mult_part_out21[238] <= P_6_5[16];
            mult_part_out21[239] <= P_2_7[37];
            mult_part_out21[240] <= P_2_7[38];
            mult_part_out21[241] <= P_5_6[12];
            mult_part_out21[242] <= P_3_7[23];
            mult_part_out21[243] <= P_9_3[18];
            mult_part_out21[244] <= P_1_8[35];
            mult_part_out21[245] <= P_8_4[13];
            mult_part_out21[246] <= P_11_1[35];
            mult_part_out21[247] <= P_4_7[11];
            mult_part_out21[248] <= P_8_3[40];
            mult_part_out21[249] <= P_1_8[40];
            mult_part_out21[250] <= P_0_10[10];
            mult_part_out21[251] <= P_2_9[1];
            mult_part_out21[252] <= P_6_6[6];
            mult_part_out21[253] <= P_11_2[18];
            mult_part_out21[254] <= P_6_6[8];
            mult_part_out21[255] <= P_9_3[30];
            mult_part_out21[256] <= P_15_0[1];
            mult_part_out21[257] <= P_10_2[39];
            mult_part_out21[258] <= P_9_3[33];
            mult_part_out21[259] <= P_3_8[16];
            mult_part_out21[260] <= P_11_3[1];
            mult_part_out21[261] <= P_0_10[21];
            mult_part_out21[262] <= P_12_2[10];
            mult_part_out21[263] <= P_4_7[27];
            mult_part_out21[264] <= P_3_8[21];
            mult_part_out21[265] <= P_5_7[12];
            mult_part_out21[266] <= P_7_6[3];
            mult_part_out21[267] <= P_10_3[25];
            mult_part_out21[268] <= P_10_4[2];
            mult_part_out21[269] <= P_1_9[36];
            mult_part_out21[270] <= P_7_5[31];
            mult_part_out21[271] <= P_8_4[39];
            mult_part_out21[272] <= P_14_1[10];
            mult_part_out21[273] <= P_14_0[35];
            mult_part_out21[274] <= P_15_0[19];
            mult_part_out21[275] <= P_4_8[15];
            mult_part_out21[276] <= P_12_3[0];
            mult_part_out21[277] <= P_1_10[20];
            mult_part_out21[278] <= P_1_10[21];
            mult_part_out21[279] <= P_1_10[22];
            mult_part_out21[280] <= P_2_9[30];
            mult_part_out21[281] <= P_7_6[18];
            mult_part_out21[282] <= P_13_2[13];
            mult_part_out21[283] <= P_15_1[4];
            mult_part_out21[284] <= P_5_7[31];
            mult_part_out21[285] <= P_13_1[40];
            mult_part_out21[286] <= P_5_8[9];
            mult_part_out21[287] <= P_3_9[20];
            mult_part_out21[288] <= P_5_8[11];
            mult_part_out21[289] <= P_2_9[39];
            mult_part_out21[290] <= P_11_3[31];
            mult_part_out21[291] <= P_7_7[4];
            mult_part_out21[292] <= P_9_5[19];
            mult_part_out21[293] <= P_12_3[17];
            mult_part_out21[294] <= P_8_5[38];
            mult_part_out21[295] <= P_14_2[9];
            mult_part_out21[296] <= P_8_6[16];
            mult_part_out21[297] <= P_6_7[27];
            mult_part_out21[298] <= P_2_10[24];
            mult_part_out21[299] <= P_3_10[8];
            mult_part_out21[300] <= P_11_4[17];
            mult_part_out21[301] <= P_11_4[18];
            mult_part_out21[302] <= P_15_1[23];
            mult_part_out21[303] <= P_11_4[20];
            mult_part_out21[304] <= P_11_4[21];
            mult_part_out21[305] <= P_8_6[25];
            mult_part_out21[306] <= P_5_9[5];

            mult_part_out22[221] <= P_0_8[29];
            mult_part_out22[222] <= P_6_5[0];
            mult_part_out22[223] <= P_10_1[29];
            mult_part_out22[224] <= P_0_9[8];
            mult_part_out22[225] <= P_6_5[3];
            mult_part_out22[226] <= P_12_0[22];
            mult_part_out22[227] <= P_2_8[1];
            mult_part_out22[228] <= P_6_4[30];
            mult_part_out22[229] <= P_9_2[28];
            mult_part_out22[230] <= P_12_0[26];
            mult_part_out22[231] <= P_11_1[20];
            mult_part_out22[232] <= P_13_0[11];
            mult_part_out22[233] <= P_13_0[12];
            mult_part_out22[234] <= P_10_2[16];
            mult_part_out22[235] <= P_5_6[6];
            mult_part_out22[236] <= P_5_6[7];
            mult_part_out22[237] <= P_5_6[8];
            mult_part_out22[238] <= P_8_4[6];
            mult_part_out22[239] <= P_2_8[13];
            mult_part_out22[240] <= P_1_9[7];
            mult_part_out22[241] <= P_9_3[16];
            mult_part_out22[242] <= P_11_2[7];
            mult_part_out22[243] <= P_0_9[27];
            mult_part_out22[244] <= P_13_0[23];
            mult_part_out22[245] <= P_0_10[5];
            mult_part_out22[246] <= P_6_5[24];
            mult_part_out22[247] <= P_13_0[26];
            mult_part_out22[248] <= P_6_5[26];
            mult_part_out22[249] <= P_13_0[28];
            mult_part_out22[250] <= P_3_7[31];
            mult_part_out22[251] <= P_13_0[30];
            mult_part_out22[252] <= P_7_4[37];
            mult_part_out22[253] <= P_1_9[20];
            mult_part_out22[254] <= P_12_1[26];
            mult_part_out22[255] <= P_1_9[22];
            mult_part_out22[256] <= P_13_1[11];
            mult_part_out22[257] <= P_3_7[38];
            mult_part_out22[258] <= P_13_0[37];
            mult_part_out22[259] <= P_9_4[10];
            mult_part_out22[260] <= P_2_8[34];
            mult_part_out22[261] <= P_2_9[11];
            mult_part_out22[262] <= P_11_2[27];
            mult_part_out22[263] <= P_5_6[34];
            mult_part_out22[264] <= P_8_5[8];
            mult_part_out22[265] <= P_1_10[8];
            mult_part_out22[266] <= P_10_4[0];
            mult_part_out22[267] <= P_15_0[12];
            mult_part_out22[268] <= P_8_4[36];
            mult_part_out22[269] <= P_8_5[13];
            mult_part_out22[270] <= P_0_10[30];
            mult_part_out22[271] <= P_8_5[15];
            mult_part_out22[272] <= P_6_7[2];
            mult_part_out22[273] <= P_11_2[38];
            mult_part_out22[274] <= P_7_6[11];
            mult_part_out22[275] <= P_15_0[20];
            mult_part_out22[276] <= P_10_3[34];
            mult_part_out22[277] <= P_14_1[15];
            mult_part_out22[278] <= P_8_5[22];
            mult_part_out22[279] <= P_14_1[17];
            mult_part_out22[280] <= P_10_3[38];
            mult_part_out22[281] <= P_8_6[1];
            mult_part_out22[282] <= P_6_7[12];
            mult_part_out22[283] <= P_8_5[27];
            mult_part_out22[284] <= P_5_8[7];
            mult_part_out22[285] <= P_6_7[15];
            mult_part_out22[286] <= P_10_4[20];
            mult_part_out22[287] <= P_4_8[27];
            mult_part_out22[288] <= P_6_7[18];
            mult_part_out22[289] <= P_5_7[36];
            mult_part_out22[290] <= P_7_6[27];
            mult_part_out22[291] <= P_12_2[39];
            mult_part_out22[292] <= P_5_8[15];
            mult_part_out22[293] <= P_15_1[14];
            mult_part_out22[294] <= P_3_9[27];
            mult_part_out22[295] <= P_7_6[32];
            mult_part_out22[296] <= P_7_6[33];
            mult_part_out22[297] <= P_10_4[31];
            mult_part_out22[298] <= P_4_9[14];
            mult_part_out22[299] <= P_15_1[20];
            mult_part_out22[300] <= P_13_2[31];
            mult_part_out22[301] <= P_7_7[14];
            mult_part_out22[302] <= P_12_4[2];
            mult_part_out22[303] <= P_14_2[17];

            mult_part_out23[238] <= P_0_9[22];
            mult_part_out23[239] <= P_6_5[17];
            mult_part_out23[240] <= P_12_0[36];
            mult_part_out23[241] <= P_2_7[39];
            mult_part_out23[242] <= P_10_3[0];
            mult_part_out23[243] <= P_4_6[31];
            mult_part_out23[244] <= P_9_3[19];
            mult_part_out23[245] <= P_13_0[24];
            mult_part_out23[246] <= P_3_7[27];
            mult_part_out23[247] <= P_13_1[2];
            mult_part_out23[248] <= P_14_0[10];
            mult_part_out23[249] <= P_0_9[33];
            mult_part_out23[250] <= P_13_0[29];
            mult_part_out23[251] <= P_2_8[25];
            mult_part_out23[252] <= P_2_8[26];
            mult_part_out23[253] <= P_10_2[35];
            mult_part_out23[254] <= P_9_4[5];
            mult_part_out23[255] <= P_11_2[20];
            mult_part_out23[256] <= P_13_0[35];
            mult_part_out23[257] <= P_9_4[8];
            mult_part_out23[258] <= P_15_0[3];
            mult_part_out23[259] <= P_7_5[20];
            mult_part_out23[260] <= P_11_2[25];
            mult_part_out23[261] <= P_15_0[6];
            mult_part_out23[262] <= P_10_3[20];
            mult_part_out23[263] <= P_4_8[3];
            mult_part_out23[264] <= P_0_10[24];
            mult_part_out23[265] <= P_4_8[5];
            mult_part_out23[266] <= P_11_3[7];
            mult_part_out23[267] <= P_5_6[38];
            mult_part_out23[268] <= P_11_2[33];
            mult_part_out23[269] <= P_3_9[2];
            mult_part_out23[270] <= P_8_4[38];
            mult_part_out23[271] <= P_13_2[2];
            mult_part_out23[272] <= P_3_9[5];
            mult_part_out23[273] <= P_13_1[28];
            mult_part_out23[274] <= P_4_8[14];
            mult_part_out23[275] <= P_4_7[39];
            mult_part_out23[276] <= P_4_8[16];
            mult_part_out23[277] <= P_5_7[24];
            mult_part_out23[278] <= P_10_3[36];
            mult_part_out23[279] <= P_12_2[27];
            mult_part_out23[280] <= P_13_2[11];
            mult_part_out23[281] <= P_12_3[5];
            mult_part_out23[282] <= P_15_1[3];
            mult_part_out23[283] <= P_1_10[26];
            mult_part_out23[284] <= P_8_6[4];
            mult_part_out23[285] <= P_2_9[35];
            mult_part_out23[286] <= P_6_6[40];
            mult_part_out23[287] <= P_5_8[10];
            mult_part_out23[288] <= P_13_2[19];
            mult_part_out23[289] <= P_8_5[33];

            mult_part_out24[240] <= P_5_6[11];
            mult_part_out24[241] <= P_8_3[33];
            mult_part_out24[242] <= P_9_3[17];
            mult_part_out24[243] <= P_5_6[14];
            mult_part_out24[244] <= P_11_1[33];
            mult_part_out24[245] <= P_1_8[36];
            mult_part_out24[246] <= P_5_6[17];
            mult_part_out24[247] <= P_12_1[19];
            mult_part_out24[248] <= P_0_9[32];
            mult_part_out24[249] <= P_14_0[11];
            mult_part_out24[250] <= P_2_9[0];
            mult_part_out24[251] <= P_6_5[29];
            mult_part_out24[252] <= P_8_4[20];
            mult_part_out24[253] <= P_6_5[31];
            mult_part_out24[254] <= P_2_8[28];
            mult_part_out24[255] <= P_0_9[39];
            mult_part_out24[256] <= P_0_10[16];
            mult_part_out24[257] <= P_1_10[0];
            mult_part_out24[258] <= P_6_6[12];
            mult_part_out24[259] <= P_12_2[7];
            mult_part_out24[260] <= P_15_0[5];
            mult_part_out24[261] <= P_1_9[28];
            mult_part_out24[262] <= P_11_3[3];
            mult_part_out24[263] <= P_9_3[38];
            mult_part_out24[264] <= P_1_9[31];
            mult_part_out24[265] <= P_6_6[19];
            mult_part_out24[266] <= P_14_1[4];
            mult_part_out24[267] <= P_3_9[0];
            mult_part_out24[268] <= P_15_0[13];
            mult_part_out24[269] <= P_11_2[34];
            mult_part_out24[270] <= P_6_7[0];
            mult_part_out24[271] <= P_6_6[25];
            mult_part_out24[272] <= P_11_3[13];
            mult_part_out24[273] <= P_10_4[7];
            mult_part_out24[274] <= P_14_1[12];
            mult_part_out24[275] <= P_11_3[16];
            mult_part_out24[276] <= P_7_6[13];
            mult_part_out24[277] <= P_10_3[35];
            mult_part_out24[278] <= P_11_3[19];
            mult_part_out24[279] <= P_13_2[10];

            mult_part_out25[255] <= P_10_2[37];
            mult_part_out25[256] <= P_1_9[23];
            mult_part_out25[257] <= P_4_7[21];
            mult_part_out25[258] <= P_5_6[29];
            mult_part_out25[259] <= P_4_7[23];
            mult_part_out25[260] <= P_6_5[38];
            mult_part_out25[261] <= P_9_3[36];
            mult_part_out25[262] <= P_14_1[0];
            mult_part_out25[263] <= P_0_10[23];
            mult_part_out25[264] <= P_11_3[5];
            mult_part_out25[265] <= P_12_1[37];
            mult_part_out25[266] <= P_14_0[28];
            mult_part_out25[267] <= P_11_2[32];
            mult_part_out25[268] <= P_7_6[5];
            mult_part_out25[269] <= P_7_6[6];
            mult_part_out25[270] <= P_7_6[7];
            mult_part_out25[271] <= P_7_5[32];
            mult_part_out25[272] <= P_8_5[16];

        end
endmodule
